PK
     �;\�	V���  ��     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_0":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_28"],"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_1":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_24"],"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_2":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_11"],"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_3":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_8"],"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_4":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6"],"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_5":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33"],"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_6":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2"],"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_7":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7"],"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_0":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_29"],"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_1":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_25"],"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_2":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_12"],"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_3":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_9"],"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_4":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6"],"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_5":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33"],"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_6":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2"],"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_7":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7"],"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_0":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_27"],"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_1":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_26"],"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_2":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_13"],"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_3":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_14"],"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_4":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6"],"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_5":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33"],"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_6":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2"],"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_7":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_0":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_1":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2":["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_6","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_6","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_6","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_6"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_3":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_4":["pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_2"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_5":["pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_3"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6":["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_4","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_4","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_4","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_4"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7":["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_7","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_7","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_7","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_7"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_8":["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_3"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_9":["pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_3"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_10":["pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_1"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_11":["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_2"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_12":["pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_2"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_13":["pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_2"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_14":["pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_3"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_15":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_16":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_17":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_18":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_19":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_20":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_21":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_22":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_23":["pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_0"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_24":["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_1"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_25":["pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_1"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_26":["pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_1"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_27":["pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_0"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_28":["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_0"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_29":["pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_0"],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_30":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_31":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_32":[],"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33":["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_5","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_5","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_5","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_5"],"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_0":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_23"],"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_1":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_10"],"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_2":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_4"],"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_3":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_5"],"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_4":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6"],"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_5":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33"],"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_6":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2"],"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_7":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7"]},"pin_to_color":{"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_0":"#9141ac","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_1":"#ff7800","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_2":"#1a5fb4","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_3":"#deddda","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_4":"#26a269","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_5":"#000000","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_6":"#e01b24","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_7":"#ffe502","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_0":"#9141ac","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_1":"#ff7800","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_2":"#1c71d8","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_3":"#deddda","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_4":"#26a269","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_5":"#000000","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_6":"#e01b24","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_7":"#ffe502","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_0":"#7544B1","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_1":"#ff7800","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_2":"#1c71d8","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_3":"#deddda","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_4":"#26a269","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_5":"#000000","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_6":"#e01b24","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_7":"#ffe502","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_0":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_1":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2":"#e01b24","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_3":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_4":"#1c71d8","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_5":"#deddda","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6":"#26a269","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7":"#ffe502","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_8":"#deddda","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_9":"#deddda","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_10":"#ff7800","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_11":"#1a5fb4","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_12":"#1c71d8","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_13":"#1c71d8","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_14":"#deddda","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_15":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_16":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_17":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_18":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_19":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_20":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_21":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_22":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_23":"#7A4782","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_24":"#ff7800","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_25":"#ff7800","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_26":"#ff7800","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_27":"#7544B1","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_28":"#9141ac","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_29":"#9141ac","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_30":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_31":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_32":"#000000","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33":"#000000","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_0":"#7A4782","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_1":"#ff7800","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_2":"#1c71d8","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_3":"#deddda","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_4":"#26a269","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_5":"#000000","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_6":"#e01b24","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_7":"#ffe502"},"pin_to_state":{"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_0":"neutral","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_1":"neutral","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_2":"neutral","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_3":"neutral","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_4":"neutral","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_5":"neutral","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_6":"neutral","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_7":"neutral","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_0":"neutral","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_1":"neutral","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_2":"neutral","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_3":"neutral","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_4":"neutral","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_5":"neutral","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_6":"neutral","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_7":"neutral","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_0":"neutral","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_1":"neutral","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_2":"neutral","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_3":"neutral","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_4":"neutral","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_5":"neutral","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_6":"neutral","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_7":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_0":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_1":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_3":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_4":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_5":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_8":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_9":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_10":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_11":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_12":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_13":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_14":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_15":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_16":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_17":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_18":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_19":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_20":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_21":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_22":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_23":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_24":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_25":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_26":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_27":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_28":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_29":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_30":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_31":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_32":"neutral","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33":"neutral","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_0":"neutral","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_1":"neutral","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_2":"neutral","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_3":"neutral","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_4":"neutral","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_5":"neutral","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_6":"neutral","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_7":"neutral"},"next_color_idx":30,"wires_placed_in_order":[["pin-type-component_9f9ee855-d43e-4d4a-adca-2df888b168e5_2","pin-type-component_eb92350a-0fcf-4f4e-96c6-d3eb2fae7b73_16"],["pin-type-component_eb92350a-0fcf-4f4e-96c6-d3eb2fae7b73_15","pin-type-component_9f9ee855-d43e-4d4a-adca-2df888b168e5_0"],["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_5","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_2"],["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_6","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_3"],["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_7","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_9"],["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_4","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_4"],["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_2","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_10"],["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_0","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_5"],["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_1","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_6"],["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_3","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_7"],["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_5","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_5"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_5"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_6"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_5"],["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_6","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_6"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_6"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_6"],["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_7","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_7"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_7"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_7"],["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_4","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_4"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_4"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_4"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_11","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_2"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_8","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_3"],["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_1","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_24"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_28","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_0"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_12","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_2"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_9","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_3"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_25","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_1"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_29","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_0"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_13","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_2"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_14","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_3"],["pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_1","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_26"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_27","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_0"],["pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_2","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_4"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_5","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_3"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_10","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_1"],["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_23","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_0"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_9f9ee855-d43e-4d4a-adca-2df888b168e5_2","pin-type-component_eb92350a-0fcf-4f4e-96c6-d3eb2fae7b73_16"]]],[[],[["pin-type-component_eb92350a-0fcf-4f4e-96c6-d3eb2fae7b73_15","pin-type-component_9f9ee855-d43e-4d4a-adca-2df888b168e5_0"]]],[[["pin-type-component_9f9ee855-d43e-4d4a-adca-2df888b168e5_0","pin-type-component_eb92350a-0fcf-4f4e-96c6-d3eb2fae7b73_15"]],[]],[[["pin-type-component_9f9ee855-d43e-4d4a-adca-2df888b168e5_2","pin-type-component_eb92350a-0fcf-4f4e-96c6-d3eb2fae7b73_16"]],[]],[[],[["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_5","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_2"]]],[[],[["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_6","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_3"]]],[[],[["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_7","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_9"]]],[[],[["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_4","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_4"]]],[[],[["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_2","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_10"]]],[[],[["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_0","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_5"]]],[[],[["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_1","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_6"]]],[[],[["pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_3","pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_7"]]],[[["pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_5","pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_0"]],[]],[[["pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_6","pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_1"]],[]],[[["pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_10","pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_2"]],[]],[[["pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_7","pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_3"]],[]],[[["pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_4","pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_4"]],[]],[[["pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_2","pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_5"]],[]],[[["pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_3","pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_6"]],[]],[[["pin-type-component_b2d27f14-8080-4f7c-ba98-af4c7a0388f1_9","pin-type-component_c21b7807-a540-4804-9031-bd43316b25cb_7"]],[]],[[],[["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_5","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_5"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_5"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_6"]]],[[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_6"]],[]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_5"]]],[[],[["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_6","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_6"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_6"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_6"]]],[[],[["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_7","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_7"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_7"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_7"]]],[[],[["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_4","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_4"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_4"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_4"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_11","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_2"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_8","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_3"]]],[[],[["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_1","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_24"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_28","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_0"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_12","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_2"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_9","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_3"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_25","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_1"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_29","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_0"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_13","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_2"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_14","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_3"]]],[[],[["pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_1","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_26"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_27","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_0"]]],[[],[["pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_2","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_4"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_5","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_3"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_10","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_1"]]],[[],[["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_23","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_0"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_0":"0000000000000007","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_1":"0000000000000006","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_2":"0000000000000004","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_3":"0000000000000005","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_4":"0000000000000003","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_5":"0000000000000000","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_6":"0000000000000001","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_7":"0000000000000002","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_0":"0000000000000011","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_1":"0000000000000010","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_2":"0000000000000008","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_3":"0000000000000009","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_4":"0000000000000003","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_5":"0000000000000000","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_6":"0000000000000001","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_7":"0000000000000002","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_0":"0000000000000015","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_1":"0000000000000014","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_2":"0000000000000012","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_3":"0000000000000013","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_4":"0000000000000003","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_5":"0000000000000000","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_6":"0000000000000001","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_7":"0000000000000002","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_0":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_1":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2":"0000000000000001","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_3":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_4":"0000000000000016","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_5":"0000000000000017","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6":"0000000000000003","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7":"0000000000000002","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_8":"0000000000000005","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_9":"0000000000000009","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_10":"0000000000000018","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_11":"0000000000000004","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_12":"0000000000000008","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_13":"0000000000000012","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_14":"0000000000000013","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_15":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_16":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_17":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_18":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_19":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_20":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_21":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_22":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_23":"0000000000000019","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_24":"0000000000000006","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_25":"0000000000000010","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_26":"0000000000000014","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_27":"0000000000000015","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_28":"0000000000000007","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_29":"0000000000000011","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_30":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_31":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_32":"_","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33":"0000000000000000","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_0":"0000000000000019","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_1":"0000000000000018","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_2":"0000000000000016","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_3":"0000000000000017","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_4":"0000000000000003","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_5":"0000000000000000","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_6":"0000000000000001","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_7":"0000000000000002"},"component_id_to_pins":{"0f06abbd-d03a-41f1-879e-bbecb11561de":["0","1","2","3","4","5","6","7"],"da03ea67-c1db-4038-9ba4-7f277a2ad54d":["0","1","2","3","4","5","6","7"],"b0c91a1d-95ba-468f-92c7-e223cc8a5a6a":["0","1","2","3","4","5","6","7"],"614f80c7-1e8b-41bd-90b7-273d7fbb8fa0":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31","32","33"],"8ccf355b-84bc-4e04-bcff-fb13ab174d6f":["0","1","2","3","4","5","6","7"],"0bcf3cd5-deb9-4ef7-9a1f-48c8812fd931":[]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_5","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_5","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_5","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_5"],"0000000000000001":["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_6","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_6","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_6","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_6"],"0000000000000002":["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_7","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_7","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_7","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_7"],"0000000000000003":["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_4","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_4","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_4","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_4"],"0000000000000004":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_11","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_2"],"0000000000000005":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_8","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_3"],"0000000000000006":["pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_1","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_24"],"0000000000000007":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_28","pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_0"],"0000000000000008":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_12","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_2"],"0000000000000009":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_9","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_3"],"0000000000000010":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_25","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_1"],"0000000000000011":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_29","pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_0"],"0000000000000012":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_13","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_2"],"0000000000000013":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_14","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_3"],"0000000000000014":["pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_1","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_26"],"0000000000000015":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_27","pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_0"],"0000000000000016":["pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_2","pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_4"],"0000000000000017":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_5","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_3"],"0000000000000018":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_10","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_1"],"0000000000000019":["pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_23","pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_0"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000007":"Net 7","0000000000000008":"Net 8","0000000000000009":"Net 9","0000000000000010":"Net 10","0000000000000011":"Net 11","0000000000000012":"Net 12","0000000000000013":"Net 13","0000000000000014":"Net 14","0000000000000015":"Net 15","0000000000000016":"Net 16","0000000000000017":"Net 17","0000000000000018":"Net 18","0000000000000019":"Net 19"},"all_breadboard_info_list":[],"breadboard_info_list":[],"componentsData":[{"compProperties":{},"position":[-81.37612550000003,97.94992550000002],"typeId":"175fa3e3-2b65-451c-aa10-715821aab4fa","componentVersion":1,"instanceId":"0f06abbd-d03a-41f1-879e-bbecb11561de","orientation":"right","circleData":[[-57.499999999999986,230],[-57.288819499999974,215.00590550000004],[-71.43818900000001,215.42826649999995],[-71.86061,230.21118050000007],[-86.009981,230.63354300000003],[-101.00407549999996,231.2671445000001],[-100.58171299999997,216.06181100000003],[-86.22116149999998,215.63944849999996]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[128.62387450000006,97.94992550000008],"typeId":"175fa3e3-2b65-451c-aa10-715821aab4fa","componentVersion":1,"instanceId":"da03ea67-c1db-4038-9ba4-7f277a2ad54d","orientation":"right","circleData":[[152.5,230],[152.7111805,215.00590550000004],[138.56181099999998,215.42826649999995],[138.13939,230.21118050000007],[123.99001900000002,230.63354300000003],[108.99592450000006,231.2671445000001],[109.41828700000002,216.06181100000003],[123.7788385,215.63944849999996]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[338.62387449999994,97.94992549999998],"typeId":"175fa3e3-2b65-451c-aa10-715821aab4fa","componentVersion":1,"instanceId":"b0c91a1d-95ba-468f-92c7-e223cc8a5a6a","orientation":"right","circleData":[[362.5,230],[362.71118049999995,215.00590550000004],[348.5618109999999,215.42826649999995],[348.13938999999993,230.21118050000007],[333.99001899999996,230.63354300000003],[318.9959245,231.2671445000001],[319.41828699999996,216.06181100000003],[333.7788384999999,215.63944849999996]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[152.2592935,544.9169675],"typeId":"b3fc962b-f486-96af-9567-1bc372583e0e","componentVersion":2,"instanceId":"614f80c7-1e8b-41bd-90b7-273d7fbb8fa0","orientation":"up","circleData":[[107.5,545.0000000000001],[122.49993850000004,545.0000000000001],[85,417.50000000000006],[85,432.50000000000006],[85,447.50000000000006],[85,462.50000000000006],[85,477.50000000000006],[85,492.50000000000006],[85,507.50000000000006],[85,522.5],[85,537.5],[85,552.5000000000001],[85,567.5000000000001],[85,582.5000000000001],[85,597.5000000000001],[85,612.5000000000001],[85,627.5000000000003],[85,642.5000000000003],[221.52100000000002,643.4345000000004],[221.52100000000002,628.4420000000003],[221.93650000000002,612.2855000000003],[220,597.5000000000001],[220,582.5000000000001],[220,567.5000000000001],[220,552.5000000000001],[220,537.5],[220,522.5],[220,507.50000000000006],[220,492.50000000000006],[220,477.50000000000006],[220,462.50000000000006],[220,447.50000000000006],[220,432.50000000000006],[220,417.50000000000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[548.6238744999999,97.94992549999999],"typeId":"175fa3e3-2b65-451c-aa10-715821aab4fa","componentVersion":1,"instanceId":"8ccf355b-84bc-4e04-bcff-fb13ab174d6f","orientation":"right","circleData":[[572.5,230],[572.7111805,215.00590549999998],[558.5618109999999,215.4282664999999],[558.1393899999999,230.21118050000007],[543.990019,230.63354300000003],[528.9959245,231.2671445000001],[529.418287,216.06181099999998],[543.7788384999999,215.6394484999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"ESP32 C6","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[152.23712517953936,503.9748794087601],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"0bcf3cd5-deb9-4ef7-9a1f-48c8812fd931","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-59.68787","left":"-185.86435","width":"838.97645","height":"786.83664","x":"-185.86435","y":"-59.68787"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_5\",\"endPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33\",\"rawStartPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_5\",\"rawEndPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-101.0040755000_231.2671445000\\\",\\\"-101.0040755000_357.5000000000\\\",\\\"242.5000000000_357.5000000000\\\",\\\"242.5000000000_417.5000000000\\\",\\\"220.0000000000_417.5000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33\",\"endPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_5\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33\",\"rawEndPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"220.0000000000_417.5000000000\\\",\\\"242.5000000000_417.5000000000\\\",\\\"242.5000000000_320.0000000000\\\",\\\"108.9959245000_320.0000000000\\\",\\\"108.9959245000_231.2671445000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33\",\"endPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_5\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33\",\"rawEndPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"220.0000000000_417.5000000000\\\",\\\"318.9959245000_417.5000000000\\\",\\\"318.9959245000_231.2671445000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33\",\"endPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_5\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_33\",\"rawEndPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"220.0000000000_417.5000000000\\\",\\\"528.9959245000_417.5000000000\\\",\\\"528.9959245000_231.2671445000\\\"]}\"}","{\"color\":\"#e01b24\",\"startPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_6\",\"endPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2\",\"rawStartPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_6\",\"rawEndPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-100.5817130000_216.0618110000\\\",\\\"-125.0000000000_216.0618110000\\\",\\\"-125.0000000000_417.5000000000\\\",\\\"85.0000000000_417.5000000000\\\"]}\"}","{\"color\":\"#e01b24\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2\",\"endPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_6\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2\",\"rawEndPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_417.5000000000\\\",\\\"55.0000000000_417.5000000000\\\",\\\"55.0000000000_216.0618110000\\\",\\\"109.4182870000_216.0618110000\\\"]}\"}","{\"color\":\"#e01b24\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2\",\"endPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_6\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2\",\"rawEndPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_417.5000000000\\\",\\\"55.0000000000_417.5000000000\\\",\\\"55.0000000000_282.5000000000\\\",\\\"257.5000000000_282.5000000000\\\",\\\"257.5000000000_216.0618110000\\\",\\\"319.4182870000_216.0618110000\\\"]}\"}","{\"color\":\"#e01b24\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2\",\"endPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_6\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_2\",\"rawEndPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_417.5000000000\\\",\\\"55.0000000000_417.5000000000\\\",\\\"55.0000000000_282.5000000000\\\",\\\"467.5000000000_282.5000000000\\\",\\\"467.5000000000_216.0618110000\\\",\\\"529.4182870000_216.0618110000\\\"]}\"}","{\"color\":\"#ffe502\",\"startPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_7\",\"endPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7\",\"rawStartPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_7\",\"rawEndPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-86.2211615000_215.6394485000\\\",\\\"-86.2211615000_200.0000000000\\\",\\\"-147.5000000000_200.0000000000\\\",\\\"-147.5000000000_492.5000000000\\\",\\\"85.0000000000_492.5000000000\\\"]}\"}","{\"color\":\"#ffe502\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7\",\"endPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_7\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7\",\"rawEndPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_492.5000000000\\\",\\\"17.5000000000_492.5000000000\\\",\\\"17.5000000000_200.0000000000\\\",\\\"123.7788385000_200.0000000000\\\",\\\"123.7788385000_215.6394485000\\\"]}\"}","{\"color\":\"#ffe502\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7\",\"endPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_7\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7\",\"rawEndPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_492.5000000000\\\",\\\"17.5000000000_492.5000000000\\\",\\\"17.5000000000_200.0000000000\\\",\\\"333.7788385000_200.0000000000\\\",\\\"333.7788385000_215.6394485000\\\"]}\"}","{\"color\":\"#ffe502\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7\",\"endPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_7\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_7\",\"rawEndPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_492.5000000000\\\",\\\"17.5000000000_492.5000000000\\\",\\\"17.5000000000_200.0000000000\\\",\\\"543.7788385000_200.0000000000\\\",\\\"543.7788385000_215.6394485000\\\"]}\"}","{\"color\":\"#26a269\",\"startPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_4\",\"endPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6\",\"rawStartPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_4\",\"rawEndPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-86.0099810000_230.6335430000\\\",\\\"-86.0099810000_477.5000000000\\\",\\\"85.0000000000_477.5000000000\\\"]}\"}","{\"color\":\"#26a269\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6\",\"endPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_4\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6\",\"rawEndPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_477.5000000000\\\",\\\"-87.5000000000_477.5000000000\\\",\\\"-87.5000000000_260.0000000000\\\",\\\"123.9900190000_260.0000000000\\\",\\\"123.9900190000_230.6335430000\\\"]}\"}","{\"color\":\"#26a269\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6\",\"endPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_4\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6\",\"rawEndPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_477.5000000000\\\",\\\"-87.5000000000_477.5000000000\\\",\\\"-87.5000000000_260.0000000000\\\",\\\"333.9900190000_260.0000000000\\\",\\\"333.9900190000_230.6335430000\\\"]}\"}","{\"color\":\"#26a269\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6\",\"endPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_4\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_6\",\"rawEndPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_477.5000000000\\\",\\\"-87.5000000000_477.5000000000\\\",\\\"-87.5000000000_260.0000000000\\\",\\\"543.9900190000_260.0000000000\\\",\\\"543.9900190000_230.6335430000\\\"]}\"}","{\"color\":\"#1a5fb4\",\"startPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_2\",\"endPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_11\",\"rawStartPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_2\",\"rawEndPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_11\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-71.4381890000_215.4282665000\\\",\\\"-71.4381890000_200.0000000000\\\",\\\"-12.5000000000_200.0000000000\\\",\\\"-12.5000000000_552.5000000000\\\",\\\"85.0000000000_552.5000000000\\\"]}\"}","{\"color\":\"#deddda\",\"startPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_3\",\"endPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_8\",\"rawStartPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_3\",\"rawEndPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_8\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-71.8606100000_230.2111805000\\\",\\\"-71.8606100000_507.5000000000\\\",\\\"85.0000000000_507.5000000000\\\"]}\"}","{\"color\":\"#ff7800\",\"startPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_1\",\"endPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_24\",\"rawStartPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_1\",\"rawEndPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_24\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-57.2888195000_215.0059055000\\\",\\\"-42.5000000000_215.0059055000\\\",\\\"-42.5000000000_740.0000000000\\\",\\\"242.5000000000_740.0000000000\\\",\\\"242.5000000000_552.5000000000\\\",\\\"220.0000000000_552.5000000000\\\"]}\"}","{\"color\":\"#9141ac\",\"startPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_0\",\"endPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_28\",\"rawStartPinId\":\"pin-type-component_0f06abbd-d03a-41f1-879e-bbecb11561de_0\",\"rawEndPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_28\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-57.5000000000_230.0000000000\\\",\\\"-57.5000000000_762.5000000000\\\",\\\"265.0000000000_762.5000000000\\\",\\\"265.0000000000_492.5000000000\\\",\\\"220.0000000000_492.5000000000\\\"]}\"}","{\"color\":\"#1c71d8\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_12\",\"endPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_2\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_12\",\"rawEndPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_567.5000000000\\\",\\\"-222.5000000000_567.5000000000\\\",\\\"-222.5000000000_177.5000000000\\\",\\\"138.5618110000_177.5000000000\\\",\\\"138.5618110000_215.4282665000\\\"]}\"}","{\"color\":\"#deddda\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_9\",\"endPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_3\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_9\",\"rawEndPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_522.5000000000\\\",\\\"-245.0000000000_522.5000000000\\\",\\\"-245.0000000000_297.5000000000\\\",\\\"138.1393900000_297.5000000000\\\",\\\"138.1393900000_230.2111805000\\\"]}\"}","{\"color\":\"#ff7800\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_25\",\"endPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_1\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_25\",\"rawEndPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"220.0000000000_537.5000000000\\\",\\\"280.0000000000_537.5000000000\\\",\\\"280.0000000000_177.5000000000\\\",\\\"152.7111805000_177.5000000000\\\",\\\"152.7111805000_215.0059055000\\\"]}\"}","{\"color\":\"#9141ac\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_29\",\"endPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_0\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_29\",\"rawEndPinId\":\"pin-type-component_da03ea67-c1db-4038-9ba4-7f277a2ad54d_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"220.0000000000_477.5000000000\\\",\\\"265.0000000000_477.5000000000\\\",\\\"265.0000000000_297.5000000000\\\",\\\"152.5000000000_297.5000000000\\\",\\\"152.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#1c71d8\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_13\",\"endPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_2\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_13\",\"rawEndPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_582.5000000000\\\",\\\"62.5000000000_582.5000000000\\\",\\\"62.5000000000_785.0000000000\\\",\\\"400.0000000000_785.0000000000\\\",\\\"400.0000000000_177.5000000000\\\",\\\"348.5618110000_177.5000000000\\\",\\\"348.5618110000_215.4282665000\\\"]}\"}","{\"color\":\"#deddda\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_14\",\"endPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_3\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_14\",\"rawEndPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_597.5000000000\\\",\\\"40.0000000000_597.5000000000\\\",\\\"40.0000000000_815.0000000000\\\",\\\"348.1393900000_815.0000000000\\\",\\\"348.1393900000_230.2111805000\\\"]}\"}","{\"color\":\"#ff7800\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_26\",\"endPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_1\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_26\",\"rawEndPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"220.0000000000_522.5000000000\\\",\\\"385.0000000000_522.5000000000\\\",\\\"385.0000000000_215.0059055000\\\",\\\"362.7111805000_215.0059055000\\\"]}\"}","{\"color\":\"#7544B1\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_27\",\"endPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_0\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_27\",\"rawEndPinId\":\"pin-type-component_b0c91a1d-95ba-468f-92c7-e223cc8a5a6a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"220.0000000000_507.5000000000\\\",\\\"362.5000000000_507.5000000000\\\",\\\"362.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#1c71d8\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_4\",\"endPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_2\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_4\",\"rawEndPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_447.5000000000\\\",\\\"32.5000000000_447.5000000000\\\",\\\"32.5000000000_155.0000000000\\\",\\\"558.5618110000_155.0000000000\\\",\\\"558.5618110000_215.4282665000\\\"]}\"}","{\"color\":\"#deddda\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_5\",\"endPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_3\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_5\",\"rawEndPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_462.5000000000\\\",\\\"2.5000000000_462.5000000000\\\",\\\"2.5000000000_837.5000000000\\\",\\\"558.1393900000_837.5000000000\\\",\\\"558.1393900000_230.2111805000\\\"]}\"}","{\"color\":\"#ff7800\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_10\",\"endPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_1\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_10\",\"rawEndPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"85.0000000000_537.5000000000\\\",\\\"17.5000000000_537.5000000000\\\",\\\"17.5000000000_860.0000000000\\\",\\\"595.0000000000_860.0000000000\\\",\\\"595.0000000000_215.0059055000\\\",\\\"572.7111805000_215.0059055000\\\"]}\"}","{\"color\":\"#7A4782\",\"startPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_23\",\"endPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_0\",\"rawStartPinId\":\"pin-type-component_614f80c7-1e8b-41bd-90b7-273d7fbb8fa0_23\",\"rawEndPinId\":\"pin-type-component_8ccf355b-84bc-4e04-bcff-fb13ab174d6f_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"220.0000000000_567.5000000000\\\",\\\"572.5000000000_567.5000000000\\\",\\\"572.5000000000_230.0000000000\\\"]}\"}"],"projectDescription":""}PK
     �;\               jsons/PK
     �;\>�a)  a)     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"WeAct 1.54 E-paper module","category":["User Defined"],"id":"175fa3e3-2b65-451c-aa10-715821aab4fa","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"f679dfe1-7b61-46f4-bc7c-d69b61239140.png","iconPic":"f78ae6cb-3b21-49f8-a0a0-4b83f9561715.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"19.68504","numDisplayRows":"12.59843","pins":[{"uniquePinIdString":"0","positionMil":"1864.58583,789.09567","isAnchorPin":true,"label":"BUSY"},{"uniquePinIdString":"1","positionMil":"1764.62520,790.50354","isAnchorPin":false,"label":"RES"},{"uniquePinIdString":"2","positionMil":"1767.44094,696.17441","isAnchorPin":false,"label":"CS"},{"uniquePinIdString":"3","positionMil":"1865.99370,693.35827","isAnchorPin":false,"label":"D/C"},{"uniquePinIdString":"4","positionMil":"1868.80945,599.02913","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"5","positionMil":"1873.03346,499.06850","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1771.66457,501.88425","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"7","positionMil":"1768.84882,597.62126","isAnchorPin":false,"label":"SDA"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"WeAct 1.54 E-paper module","category":["User Defined"],"id":"175fa3e3-2b65-451c-aa10-715821aab4fa","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"f679dfe1-7b61-46f4-bc7c-d69b61239140.png","iconPic":"f78ae6cb-3b21-49f8-a0a0-4b83f9561715.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"19.68504","numDisplayRows":"12.59843","pins":[{"uniquePinIdString":"0","positionMil":"1864.58583,789.09567","isAnchorPin":true,"label":"BUSY"},{"uniquePinIdString":"1","positionMil":"1764.62520,790.50354","isAnchorPin":false,"label":"RES"},{"uniquePinIdString":"2","positionMil":"1767.44094,696.17441","isAnchorPin":false,"label":"CS"},{"uniquePinIdString":"3","positionMil":"1865.99370,693.35827","isAnchorPin":false,"label":"D/C"},{"uniquePinIdString":"4","positionMil":"1868.80945,599.02913","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"5","positionMil":"1873.03346,499.06850","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1771.66457,501.88425","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"7","positionMil":"1768.84882,597.62126","isAnchorPin":false,"label":"SDA"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"WeAct 1.54 E-paper module","category":["User Defined"],"id":"175fa3e3-2b65-451c-aa10-715821aab4fa","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"f679dfe1-7b61-46f4-bc7c-d69b61239140.png","iconPic":"f78ae6cb-3b21-49f8-a0a0-4b83f9561715.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"19.68504","numDisplayRows":"12.59843","pins":[{"uniquePinIdString":"0","positionMil":"1864.58583,789.09567","isAnchorPin":true,"label":"BUSY"},{"uniquePinIdString":"1","positionMil":"1764.62520,790.50354","isAnchorPin":false,"label":"RES"},{"uniquePinIdString":"2","positionMil":"1767.44094,696.17441","isAnchorPin":false,"label":"CS"},{"uniquePinIdString":"3","positionMil":"1865.99370,693.35827","isAnchorPin":false,"label":"D/C"},{"uniquePinIdString":"4","positionMil":"1868.80945,599.02913","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"5","positionMil":"1873.03346,499.06850","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1771.66457,501.88425","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"7","positionMil":"1768.84882,597.62126","isAnchorPin":false,"label":"SDA"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"ESP32 C6 DEVKITC 1","category":["User Defined"],"userDefined":true,"id":"b3fc962b-f486-96af-9567-1bc372583e0e","subtypeDescription":"","subtypePic":"47e6ec23-9fd2-4f79-b93f-ab3ba2a25103.png","iconPic":"5119bd54-fe8a-4b53-af25-af94989a1f77.png","imageLocation":"local_cache","componentVersion":2,"pinInfo":{"numDisplayCols":"10.00000","numDisplayRows":"22.96424","pins":[{"uniquePinIdString":"0","positionMil":"201.60471,1147.65845","isAnchorPin":true,"label":"Pin 33"},{"uniquePinIdString":"1","positionMil":"301.60430,1147.65845","isAnchorPin":false,"label":"Pin 34"},{"uniquePinIdString":"2","positionMil":"51.60471,1997.65845","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"3","positionMil":"51.60471,1897.65845","isAnchorPin":false,"label":"RST"},{"uniquePinIdString":"4","positionMil":"51.60471,1797.65845","isAnchorPin":false,"label":"GPIO 4"},{"uniquePinIdString":"5","positionMil":"51.60471,1697.65845","isAnchorPin":false,"label":"GPIO 5"},{"uniquePinIdString":"6","positionMil":"51.60471,1597.65845","isAnchorPin":false,"label":"GPIO 6"},{"uniquePinIdString":"7","positionMil":"51.60471,1497.65845","isAnchorPin":false,"label":"GPIO 7"},{"uniquePinIdString":"8","positionMil":"51.60471,1397.65845","isAnchorPin":false,"label":"GPIO 0"},{"uniquePinIdString":"9","positionMil":"51.60471,1297.65845","isAnchorPin":false,"label":"GPIO 1"},{"uniquePinIdString":"10","positionMil":"51.60471,1197.65845","isAnchorPin":false,"label":"GPIO 8"},{"uniquePinIdString":"11","positionMil":"51.60471,1097.65845","isAnchorPin":false,"label":"GPIO 10"},{"uniquePinIdString":"12","positionMil":"51.60471,997.65845","isAnchorPin":false,"label":"GPIO 11"},{"uniquePinIdString":"13","positionMil":"51.60471,897.65845","isAnchorPin":false,"label":"GPIO 2"},{"uniquePinIdString":"14","positionMil":"51.60471,797.65845","isAnchorPin":false,"label":"GPIO 3"},{"uniquePinIdString":"15","positionMil":"51.60471,697.65845","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"16","positionMil":"51.60471,597.65845","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"17","positionMil":"51.60471,497.65845","isAnchorPin":false,"label":"NC"},{"uniquePinIdString":"18","positionMil":"961.74471,491.42845","isAnchorPin":false,"label":"NC"},{"uniquePinIdString":"19","positionMil":"961.74471,591.37845","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"20","positionMil":"964.51471,699.08845","isAnchorPin":false,"label":"GPIO 12"},{"uniquePinIdString":"21","positionMil":"951.60471,797.65845","isAnchorPin":false,"label":"GPIO 13"},{"uniquePinIdString":"22","positionMil":"951.60471,897.65845","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"23","positionMil":"951.60471,997.65845","isAnchorPin":false,"label":"GPIO 9"},{"uniquePinIdString":"24","positionMil":"951.60471,1097.65845","isAnchorPin":false,"label":"GPIO 10"},{"uniquePinIdString":"25","positionMil":"951.60471,1197.65845","isAnchorPin":false,"label":"GPIO 19"},{"uniquePinIdString":"26","positionMil":"951.60471,1297.65845","isAnchorPin":false,"label":"GPIO 20"},{"uniquePinIdString":"27","positionMil":"951.60471,1397.65845","isAnchorPin":false,"label":"GPIO 21"},{"uniquePinIdString":"28","positionMil":"951.60471,1497.65845","isAnchorPin":false,"label":"GPIO 22"},{"uniquePinIdString":"29","positionMil":"951.60471,1597.65845","isAnchorPin":false,"label":"GPIO 23"},{"uniquePinIdString":"30","positionMil":"951.60471,1697.65845","isAnchorPin":false,"label":"GPIO 15"},{"uniquePinIdString":"31","positionMil":"951.60471,1797.65845","isAnchorPin":false,"label":"RX"},{"uniquePinIdString":"32","positionMil":"951.60471,1897.65845","isAnchorPin":false,"label":"TX"},{"uniquePinIdString":"33","positionMil":"951.60471,1997.65845","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"WeAct 1.54 E-paper module","category":["User Defined"],"id":"175fa3e3-2b65-451c-aa10-715821aab4fa","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"f679dfe1-7b61-46f4-bc7c-d69b61239140.png","iconPic":"f78ae6cb-3b21-49f8-a0a0-4b83f9561715.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"19.68504","numDisplayRows":"12.59843","pins":[{"uniquePinIdString":"0","positionMil":"1864.58583,789.09567","isAnchorPin":true,"label":"BUSY"},{"uniquePinIdString":"1","positionMil":"1764.62520,790.50354","isAnchorPin":false,"label":"RES"},{"uniquePinIdString":"2","positionMil":"1767.44094,696.17441","isAnchorPin":false,"label":"CS"},{"uniquePinIdString":"3","positionMil":"1865.99370,693.35827","isAnchorPin":false,"label":"D/C"},{"uniquePinIdString":"4","positionMil":"1868.80945,599.02913","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"5","positionMil":"1873.03346,499.06850","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1771.66457,501.88425","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"7","positionMil":"1768.84882,597.62126","isAnchorPin":false,"label":"SDA"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     �;\               images/PK
     �;\<jݍ�� �� /   images/f679dfe1-7b61-46f4-bc7c-d69b61239140.png�PNG

   IHDR  �  3   �5�   	pHYs  �  ��+  ��IDATx���i�eeu6|��g��gP�p�T��[��Rf�Kex+�J~��ˏ�J~�������T�e��51Ā� B Ad�hzzz�g>g����u��:�<M�wK��9g�{�ú�5���1��.|�e�}ƿ����"/b]㛼(�C��(���ʲl����v�����o2wO�g]��7�s~�����]G����{���;�_�t��Zw͢c�N�:}zO����!�f<��{����B��������s,y���Z�j������[8v�ǝhu��՛6m���:y������ښ5k�l�����s�}�嗏=�V���S�'���t8F�h||������+V���Y�ȅԲ6�����3'�&��knn]B��%>�A���v���l�O���4�Ƥ�K�w˖-��独�p������+|l����.k����?����F��ͨ˨��g��͒���y�@8��=?RO��+�Gf��nǑ�����7�v�F���`�@T�#bUc>�T�)ٚ'ۼ�j#����x����p�x��_qf���ʂ��X�Y6zV�S�EY�	(�/��ܓ�f���9�����M�}&aآ���,�\���a��A333�;���~r�B���f���͸	N#P������/�zd��<��E�O�Q1�x9�e��	�Ѯ]��iW�\�����Ov�[�h�F�<��Ɖ��WB����%>�Kx�ĉ ��+�Zx��#��'�
fw���U�6�	�ȧJ�؍Dmr�dԵ��ڠ��q?� +����K ��`�ᥘ���ڷoZ8x� �#��x>��B'q'��f�N�`ANj��q��}�Cұw��n[��899�v�'�t�_�y�:֓K6C_b�ٔ�>N��g�xv�����F5i�g?+�Z n���ѵ��}C�4���M��&yzz+�⯜,DBI��yC."��lAF=^R���=$�)l%�Ƶq�FNo�Vs�lߌM�cr0��9�5ւ!P�e5t3��g����_�O�Ѱ�Mr3�h���#�	w"�M�]�4��O����v�=~�V!�p�F�:E�� ?sBl��;��:�������_)@�X�7�v�믿�6�=D(
:�v����ggO{�!x[��hp\.iA��b@��E���KPѺu�o�~��g�3��#��Qῃ�g�kBXT��(t��/|�{�{��'1)$w�狛����<� �����f��H��9���b�?���}�C��	/�X;x�s�e#Sz5@����mh%�My��b��r��ҽ4:�㬳��#�o��E�]t���>�pTR0�� ����Ӏ>���l$�z��r��-��@!N�
�$t#�Lt.��I������<^�p}?mN+��gc?�mO�F��_�0�a��<9�\6�-��~�,���:c��v?�ֽ0̴@�A�K�l?��Q��^�޻��Y� ��TEٝ�`�c���H
��e���K�=u���b����U`Æ���ss6�2.k,*�U�=PRk)�dB<w.�7�a@��Tt��I<�/��MI\`�	Ae��T
n�^�ZP�)�Ԇ�قTd4֑E�x}�E\{�;w��ꫧ�Vm<yx�x��x�`�B�޽{�}����<���=�h�&����$�ն�(��rr���2cy ���vi"0�5B$��E���y���,����s���g��&*6�'{ۼ�(�WhӦM�.\x����ܽ�i��f[V>5��>���7�:i��B$�T��آ��-%4N����8�� ��!����P���_{)E{���A�fóy~��@�5�%��q�wZ;&��g�3\�!&��^��ejjveֈ�j�*x����b!�,6od��@\��i��7,j���FH��F� g ����oٲ��� ��(�f�5�����N>��l����_�'
�@j�0��|�;џ]�vQ"��#����.R�3�빣1E�"�N�+Hѭ�y��F?��#?��W\�����n��+V�
�B�_�Έ��7�$p�(���~��_���ha�+������)������?6�����d�;� �E��ۖ��A�)|{t����.]��j}u���ɱ1�[�j������`�q��d���d�\�L96�rIaT�V�Z��5k�Ӌ!��)�y�0�&��M�l�E��Σ3�L|�U�-aJ���o9(�ZW̸�9����j3:����$q$K��ߨ�Є8��F��Z�y-<bΪm�9i���jʆ����F�a1ٓ�A����'�����:9N���AU�f}Ux�!�B.�7���ǣ
��L�)���l����pO��`F���{��g�P����/ǯ4����q�8�Q-�����F�k�.h.���T�)B��(���<>�r������c��f,4�ȃ�oܖ��0����;+J.D�X�ʢ�u��C��F�T�9b�'w$1gI4�G�@�W^{�����o��vt��U�wL���M%}h�������SYp뚯�8:en�f �׃mj��	ͪ��lO��3��4i� �2�6����ר�&&&�9-�B��:S��4�N�E*�\��n&^���i�	���5�`W�쟁�.S�[Yw��r�|�Lc-*'��)��hh��}���<p�i�C�g�C_m�K�g��	�7�5��U�(��n���D�ˬ7� e������=(�W�#5��MW�C#PK04�hӜ�����3�vf=��4��P՚����9ӟ��31��ab�ɹ$���>c��S�v������^��L����"{�3���{�=-J�ME��-�7.���LȠ�`��<ϗ����I�4fi 1�,�9��]��3�,�ܳg4��Ʉ�Z�̭}$����"V��C�D�;��kNny۰D����O< ſ��;�s����/}�k��m���k�'r���Oh:Y^�i�Y6��{K�N ��%�/�"dʱsz�0��V�?ӻ� zl	�76_ܷ�KI�`��b�ɽ���,o6iel�0AQ�SO�ZZ\�Zfͺt��k���`|��|�V��ϩ�y�DK�.ىp����Z3��}i�ԡCs�
q����|Ac�L{��ٲ�����G������(#0��Ӡ��Q���h�h�2�2#Ct*�Ap݆v��B�=��ۮ������Z���
Ώu�H�/��8J���ѿnn~�w}��2��ȧ	^F羫�T��᪑ 9��~~a�/}�L@&6����݄�Y��*(x2k�,QRؚ���S:�����;A�D���Ƶ��e>5�%T�B�oj1�q>���ju�.�?�
A�r���F���eg�;VF�с��9�&��|���Q�^�Fʕ�(L��vُU���~�P�	ey�ቕ+����8��_�N.�c�Ax��P1|q�=��:u�w�w���z�%����ٯ����������!`v�nd������i�zժU�W���a[�����bzf�m��0�\6 �x�>h� $�N�A��>��(���D�E���X�3XQ�u�w{p!��1��I��I��$Yc�4�Dg�(5~�� ;���枅��"	����`��l���I3{BP)���RMH!Ҽ�0�0��Z$df������J�����'����1{�L��7nm���l���5��͗����.S+����}���M;�2��������l�&��i�g�^���5��l��P�מ���j�a[��d�|=�7��3���5�'�D�� S�y�L�Q�'��� N����F� ��O��71陃��c������Ӝv���$�Fp���`���L�"�J��֭?��֟�.��T����}�С���#���F�?��nݺg�}���������[o�))��^���y����7�'�:MS�Hіiށ��֭���K���'O9r$1���N6Fɢu(i^H!�i�I6�"�Ti �аwR˲}��jF(�8�)���*�?��f���&/�^M�0
���cX�DW�r��%.4��KmAc*�^�)ȧ������OR��e���y��	2�;ݒ$X膲�KN��-V�~2���Ce<��(� �Opc��������2�
luv+}N��z�.�<�@�/G�
������XE6��l�-���x�3���
dAmM�|F�.�O��c!ySTrH�I8+�_�`��&�R��N��u� ��o��Q�N���n��!Ϙ���r�N���)�����G���[��)�:�VT3��N� �B�B¢���Q&��h�A���p.SH����r�C�M����	|���q>�L:���!�8�(�R����V5�3*.u/诼��۷ONv7m�ľ�/����n'e$lٰ`x�p�ݻ�@�]�j�pݗ-�5.��^�җ���}�#���fY_��z'�!�B��D���N�8�~���.�l�ڵ�1 ��cǒrl��/�d1�"ٕ���rq-E{J��߫����3�%�qZ�+j��&��k�i(�"���w��F�g��|���Mz�9:�q{#q���};a ������ZrATߠ��^k5M�� �`/�{Z��u^��e{p/<
��È��Z�e��޷���5۷gz0�+8����o��������o=�{b�TC��k���V�N����'�ܙ�K���䨥h�����@��FO�~B�F��7,�8������ `ff�.0�l,j('�i�C�7	tT0��_�ַ���� fgO>��ӳ����ڛǲX�Ŷ�r%���۶mK�c�|��a�!P[��+���/~��Gg>����D�4z��?M9%�<�����O�t��Q ?���n��S'fo�ᆝ;w���_�=�� �؃ �4����r�������۶n|<p�얝�kr̂��$�w�$�m{??�.j�:,�u.^���CI��5p�v��И$&A�魵��'gȆP��Fd�z�s��۽a�]4J���vf�1�M3z�����2������W�%[�-��w�8Sޥ��3S��(�Z�㑞rZWk}���V�=n���u~�-��� s0��G�b��r9�l��7�n�n(eC�m��&Y���$_�҇�s��W�c�"��\f�l^�Ne�(zw&�)�,dFc4f�CR��&'���0���:�Yfͨ=7�F�z��<����W���7߼e�����{^�S�wrr..ͧP���7K"~��G��fOy�f��K/�d��-�O�8�f�SQ!Ӓ�o߾���^�nݻ��.��Z;�_e����w��/����6D̈⨙�����n��ꫯ:pprr-��)���)H�Ɇ�5Y�ɒ�縧��Y�f=$�Ǜ�Zi�WM�r�<>�QR>��д�q�
)S���o��
��2u����(�&����4Di�@��Q��bi/u�04�3=>��~���$��=�r��L��=�g�4�Rt�U�[�Բ��,�g��������u��L�����,���7�Fm�muo8��r|�����n٫���-�Liˍ����`�B;�`k���ñ���?ھ�1��i����t ���c���B2E��rBw����d=>>�}�v4������ɩ1�@-��� �B�C.�ms)����@�f͚�q��n _t�%�7o>y�4�Y�� &K@��k׾��kw�y�;.��ʥ��aM%��Et�{��я~4)̊�)]��9[סs�?�"�}���ѡ � >�v���]�L�/�!�����ڵ�6l�81����çN�$�a��^U�p�N��u7s���%�8,,���tzr��&C�����`��(0��\j��J>�Ԍ�ꂶ��wҿ2#L�[qx'�)�Ri�d�΋~o�4���5� � �)53�j�Ҍ=��N��$8&���?��n`�4&�EN�]a:K�n���V�O�[R�ik��p�8DA�im{�V<����b������s��dd?��5�w�Z�r�Q��[���B����"�Sb+��~f�6�j�{��,ѱ����u�;�)��F���|V�������)����aSDwTeH�Ah�59�_��+��/��oD�M�+'�x��]/�ٴy0�ս����..��<3����'�%�fq:��H�'��:]�ۘ�����Ǐ�\9e�Z.��㩧�z��޲e�j��� 6��$�k �k��@����'Ob�V����fo�����XO9����'N8pPrU7��wj�l�����#����F�\!������3Wy��C��[!ڔ�K�q�6ՠ��5��h��,�� ,���ɵ�eL# hd:Jp-Cs�2>Z෍w��fm�����&����f�xP�����������e��g�#9"ia�M����~لDg��_�`AD-Cʲ�Gl�~}����������c�4����Wۤ�����u���et�<9��)\�^����ga�M��;Ȃ�F	�0׎m|O��Aج56&+�A6��;6�܃��F{)+p���5����I\�z&�����Y4q���c��	�p �hc�� �u����k���F��#y���{�00���/C�'���� �K����?���>���{��\����s���]p����M�,�T�i=q�P����xd�K� �7o9X� �+�؇d�)�<�npu��n�d�F5Ph)ܣ�-jvF�
 0���KԚ�.��+��L���Xa�~�5{�u8�A(+�ٟTέV�?��0r˰���M
9��� ��[Ҽ��DFMߨ���v=�*R�߇�E�aîT�:������/~�,.��5
[����@��/����"E�Y��e^�@�X�3��Sv�T{�e�u���P!�0���e��������F�E�N���a�l���Y!�<�l�P���j�5�cd�G?���ؘ�F���I��be�)!2e����xVG���m͆��aݺ�G_C�~��7�?������yl���[7��]��+�(�$#ܣ�����Cl<p�`�|��}�N;WM�̟Z�]"���C@d��K/��裏^y��5,��HݵƊU�~�i<�@����� �q�|�ݻw߾}��o޸	�᪫�ڶm�Yg�����f�$&$ٝ�J�޽�gO���ضo��>t�ЪU+c��X��;��'�x�5{�͸ڹ�Rl%|�f$���HC��>x����72Ɯ�L��b�ق����E>�z�i��O�5.i�ä�\#���F7����V�t�0�g&��+���,����(�Xʜ�zs9p��� Y�̂�f'���lc�#)0� �����~�u~��U���$ �� �#3�^����0Δ��L-���|�т���ʫpM����ਟ|Xo�o}�\|6��ڝ�Vd�4q18;��:�7���ރۼ�i,\~���~�&�X���a�n��A7N�E�Z�K\�(�=r�0`p������oy��������zT�L���-��� �>���=��SO=�ځ���!�����A�8.�"�'N���������[���jכ0�^��ǟصkO*gʙ�E�O�_w��'�{s�6�������Бi	j�[�"�z���r��.��򍛶 �O�.��=ޯ%n���-sFC�oٹ���/^����kW��Z�0�>�ä$������vHXɠ�95֯Y�% 25k�Z
��΄�y������*������XQt�*�elvvv�(30�Ņ8nfE���SR[5���s�9�ټy#>�bl;V�trrܱ�~Ԛݒ����d�/L���a~M�ŭ���Q|�>�π��y�?������R���v�RpN��q�����X�a�]�JE-H�5E��3`>�L�D�B�k�,͸�����A0.._P�	V���yNʖe���x��� -��+�$�gv!q�23hN<������(��Ņ#�Dk��֬M����4.
k*�Z;�����d�f��W��L�p`��J,l���enq��q��tA�;��~
ͅ	Z�x�~�z�q1�d���17�k*�Y�KЫS�b`@q��2c�.���"2�m!ZHݝ�TJ�gV��VӸQ�R<Lc��Vբ�םuֺ��ȱi0��������믿~��P�a�Q��sw\p���|�#��w���;߳���Bށ��_�u��&/��Q�2��K/|�{��q��&��L4x]j����yiX��NV�q�Ds��~o3ȕ������q뭷nܰ�q��1��4���D��n$�=�E�_|�;X���I�|�����$h����3��\I�_M������t�Y�#�!�>pK����B9;��Gu?e�
�M%��g�O��ug9r����t�b�0d�(J�o��z=�@<��j�BCQ+�׵V��*�s�3����.D$hT�~�L��U�1�e�>`bԫW����R�?��7~���P6ʏ-C�wr��kG�}{�*8��Ќ�̕n�e����2	�p2?S*M1e��02gȴ�S3�ZaX�O���h�&AZ ��"�)��H�:$'K�ndd�>
�6gZT	���lܖ�SW���ӬNS����A��hW  c08{�7���ΩW�t�E�5Ha �1���l�@��"��d��1f�瀌@(�����g>���]�������F֭['b��qjw��aEڭ��a������疏|�#\x�ѣG��F��t�Xe3�K�.  �UW]��o~���������!ec8�����Q�\��x��^s�5A؞�37xm�8t�==;{:�����u�z̧ĺ�g�+���$���=	��Ї>t���NEʱ�Xe�)(ѓ:A*2�)n9��Ǎt�7@mȘ\�����JL/�2����˶����u8ʟ�K-�\Ĵ�EdXw��#�,�Ͳǰ0o�2 ��w�6�)n-�i||Rj��U���VE!��G�&�Xv����#*�=�Iql .�r��0Z-J-ĐG���ZT��\�����RرWdΐ�!s��W�S��;r����$ʆ�t���B+R$AC���"�j�b�漙(m%���%f�x��Z$�Hdpo�c�L�k��e�ZO�VB��"c3u���@ �k��R�/4{��f�<���+-��F8?��~�)�
�O��VB$�b��c7{,+y2o(�r� �ʁ>j�"d�ܖYn�TJ�l���
�s�iɪZ;@ϛy�39�i�ոm�޽ ���Xt:�����$��,&e*�a���#h�.��R
� ���O|��~�0��'��D�Tg��"/j�2�}��ʡ%�y�����@�/~�v�Z�~D�S'glu��F��e#L@bg��+=�Q"e�Ԋ={��E��1g�y@�ƍgff�Q1'gR,�>��~���I��[�FV
o��őS�a�u��EֈA�۶mÿ���ׂ��L9e����Q�K����𨵨�j��	�A��ɝ��xmG��C2���W�� �����K���=��bl��\�J�B��R1jPf��A��I�-��J�o�<��ab+�[9@�yYY���h����λ1i���k<T�1],a(��4	�ֈ����\녚�Գ�);L ��ul}�bL�Poͧ�=���x]iW�Q�ٰ})j�CK�����ݢ;�ïi�V��}6o�	��9؟��As�`Q|YD�=�O�+{����L��[ʆ�'1�a"'�3(��4W�Rf']q��*A#6l����zlp���+f�7�N�'�Z�e]�v���C`z~�w ��3��>�Ǉ��$);L�N��$=��_�U|����=��*8na�����v��Ço߾#�\�H������G�N���`��Y�Ç�^��;x�uL��bz͛���w��=�������I�6}<�xCn`��_rB�Ġt�\�H��=�.j7q��k���}����n�W~Y�e�oЍD{A|ͪ��K��x��ׅ���\�U�XL]wR>�Z�l#yU*H�[�#s�A4RktQ�O��Z��f&a�Fg����=&N�Z�*^d��)ף�X�%���¯ͪm�%�k5&b�(+�@d�U]0>G%�8ba��}��l6�Z1ؚ͝O�13���g�õ�5�eL�@��<,�m	�=[j��\���QV;��*w�#����s*r-b�HEvh�_
��B��i�lUW��dQ)�q����9Ս�)���9���rDtM��*�R���:+E��D0�	�笳�Z���ϊ;:}�D����5��$��0D��Qt@!���*<r��k�_���n���6i36�� �R�/�z�
����%�.�m��铟ڻk�#����J����p�4
�g��#���sn=��+�!��7�;��4�Bg)!��.C_���������h��a��j
C�$>���԰�<����{�(\k���w�ӘZ��e��J�EW�xa�q�J��c�X
I~�4�F��anݺOA�2Q��;c���	��8��m�&� h����a��~��&��gi�a��O��Iw���6��� C.^���ˣ�t��X�~`��k�S(W��l.5�a-j�V7i��4d4
�NT��BOq�	̆�#w�]E{�Ը�ч�d���*��5d����` �i��9�:f�6��WG
W?�v�r��0v�L[��y�:���<0B3�PUZ��f�d��Mk�u���e�D!q�8�k)-1�r�aD)�]L�Q2���ʹ/e�8�X6p�4	\X�r�w����Ve��m�쾽%�D�D���n�\�B������K/�8qb��Ր��ǻA�=��t��σR�n��دMATN��T����T���t�'���'c��Y�eW_}�\@��'V]RG�ǚ��̩N6���v%:țb���sv҄�h�S��A�opKD&�$e�R�Z�+fI,����6�/@=IY�C����<�;�e�a.Mh��v����t~���m;�\G�OE��F''Vtʱ�NJ���TJ}�Bz3����b*�3nn����6��zX����YA�\��;l��L>��|"s��Z:��2vm�@ _��L��j��������ٲ���.�����H4FeZ�cY���m�+G���	 ��Y��7�M�P��Z=
�F��$��ӣaF	��Sy�e��:>M��N��!�Ƌ�J�d�:����Y5rJo�
	u���3��l�U)��.BcMJ��4)0A�hߠ�2����==D��Ipɖ��4o2��Y�<-�<�&� �a�5хzp��`3�(Z�|��6l Բ�Y?/�F��(��b,ٳer�5l[f-����@6;���s��'�x��p��p�W�:�A�p�*|,.u�2篖�I�F���7��;Rhy�ʕ7�t���3��t��n�1����R*���,[L2�
�K1�Y�3������I���Ͷn͆�Cței��	k�WP,8� QS��A%f+Ūc`6n܈ᶴ�(>c~��������Zi1elN��C\��a��Pj��:Ӻ�l����\+�θ�$�¨X���Ur=�x�H40CB+)�s�g��R��� '��0�\�S�݊~�%��$sFt��H)��^�s�l���ka������l�4K�i���W�[Oӑ+=Ռ�L 6z`��Օ��S�#�A�◹F�����0'���I3�f\Ө�d#cQ�Ҿ땹�Ԅr��a�L��5"Q���-�!��2Eji(�mO��Fޙ��I3-�g�q0?Q���¿�!ue�=v�O�N�M�`�J6�j�&�"4#��{�7�޽���Y@d?�3ѕC�295P�G�dw�5��jBG{r��ԒEi6块����_x޹ȗR��5�vOn?����b�hI�ixt=�P��Ղ3�w��䍉ld.R[o��v�{�J�!N����1�hI��36mڴc�hLX�2Ԝ��Y���+ k������s����=h�9�@s���#�P݌�&�6�I�3�<_vD==��o������+Y)�0�3r=h��cD闀�P����,��I�%1��-Q���5�F�V?z\��C�������Y��B�ITv�B�x	/m�Z?9չ�n�:Ό(k��{�3+P�g�Uz$����Yـ;�pM�@@ɤ�MZ� eZA{6?�s�FTQYt�4�d�Ņ�!2��zn� @��.�+(��y�K�a[,Qw,I���+I$̓��aN�8#ތ�I|�3ڹ
?�EÂ g7 �T[$K��b
�ڎ �a���ab�LU�(�Ώ�_���f���¬-Jt�3j��ȥ"�lݺ���:�)
&K�O�Y+s
��-ŉh�(֘���M�P׾�-O=�����72l���=b��t�^�7��r�"%�`�l�YkD0�h|j��o~3f3�-
k퐲��F?;�+���P��d��F�5Ggylϸ^�?=��F�*���5N�:�k�֭#��(���l�����]l�W^y��6�	Z�H�щ�� ^��d#4�u�x��:B��B>��a�)��\�uf���(���槂�O����38d*�R���������&r��l\b���	`��\�t��dS,�f���G���3 ��ˤV;i�5X��,�������i]Ʈ���Z�5L��i7��k��L� &��֘�P���Fx�ƿ���^t�:zvWt��'�AلgQ-�*�^��������)���U��{��I��O19������$��wh��5x����o~���j&f����q,�^h�I��D���<��b�31_� R=hDU;:E�W�}����W�!3�a�2��s�yvk���K+��a����sY �l�=j��-Va����4�R�-�ma!���S��n�I�d��V�Xy�%�b���!���Uk�l�:�A�|P��H3�LE�dj��Ha��	���Ρ�1�r�KSU����J0���!P��{�[���z33K�/��6`�7��������@:�~+r��mW�\	pam,<� m0pS�l�����;?����8�)s5EhE���)�2�oѤnc�U��ܡSA͗�&~�¥r�v�9�kf�L���|
zŜ��ӡTC� /'d/�W������h�R!炇�B:� ��) K�)z�2����X70���Bg<�G�4�ER7\J='�W�x�/-���ć:�����d�-�R�(f����>��T�/�b3DOx�\�VaN*%���@%��31u/�v�Y)�H�9Err�B��k���`�,w�<���<�^BT�q\f�W1��J!ʒ�pݗ��)æ9;���,��a����m�-���{i�;y�-żX�RK�$�v���#9n��-�5�ʤa��>^�'�m:(6�����ݜ�G��l�B��w�1�� �ռV��M�i���Bw	c��į�kכ�KΉ5�}�r��T�fcQFb$�4�v�Z��bo)��'6�_#Χ���hps�����a
����,`߾}�9L�N� �Q�A�<ڜN$>nZ^\,��#�x��I[-��u�p��eO�n�	��M�S���r����S����_�3 (�^���y�{�޼�J(��������Ϟ=~����!Cʦ�ĳ�Ix~bDj�c���\�̓	ɚ��L���"Yh���rO��jr�fP��5Z���Rh6]�=%/:�yB�ٯ�d����L��	��*R\ԡ���}�eǎ��Z��21�$YQ�v�R���$�ܟ���1F�H)�p��څ�����̩tQ��9��]X��|;_����o�ꪫ�%C�>�sj���:�	�х�s�����l���ȧ0mf�(���� �epLWCf�`�썶4�� Ld�)o�Ƞ_��9h�%��v2���Q/���H��t�#�Z������~�{�m1|�v�ȣ��|=���9�$�\�uB�]�c�o�%Ũ�c2Ћ�n5�Iu��R�c���r��`F_k
��$A'N������s,�,߁�M`����o;wlb7Ċ���I��p%��Ǔ�IV�y���@64i1j��\̂�gg ;q-m)Z�u����W�x�'q����H�k�3R��1/T+]E VZ���&&�Z����÷�r˭���� 8��I9�m�Y���[�l�ַ�5U�����'S�s�΁� u�j����E░���kH�Ừј�t�S}�^�7Rp-~K�=��Y�r%�������.{����ѓ낂H�g���Y�dLU軃��d�?������ ����9�[�l�ڸq��E	)N��F���_|�_�����o��F�#��CO�_��7v�1�:Y��b�+�q����o&e3��P!������Ȓ0,=$7�_ГR�C�{KW�LzIbM8�>�.ʤ��S�>�܏�}�;�ٺu�W^-U���D=*3��+���҆�r��o�ۜ��X��7mѷȲ�I@�L�&����x,g:F&�+-������H�A}9�L�%H��i�)�D>$�Q��b���A�sL��.����;6�I捈�������9X@��Cރ��D�R��l�e@�V����a���/!���J9S�}�M��Z��̣k�-��2�Y�R�?;th�Y8_qpPz0(ʆ�Z������45����TJ:<mVo.n.y��^v #B��:�kg�|��B���Ϟ<]p�9+��v�N��>���ڼ(�vfDJ�A�Iv�R��ݛrg�VT���QY�x��M�d�����o!^|3����FL$�������ٸ袋���wNMMI�q�b�Qȼ_w�u����c�>���YV�d��\�fMnA*3PȪ�x�4:��x�mh�m�FF��A�T��L�|���?����w�}P��tj-:a����b Ai��7LF�(��.�-V��H0BO�*��g�ͧ��$?���?��Ͽ������}ӛ�D��[�̒�3�~6�7@�{��'Y��?==�{�oߎ��WL�5�\ e*]�r\ðXm���S��[���AJ'� aA�+�b�.Pci����S�l�F�` �eM��s����,�/jR;�@-e�k#��zGw�
��dtJg�8�R�&���ZA������W�/.�M�N皚�TA!i�n Ε��jr��l�R� �cbl�/�҃8U�t�x�X�	�wjȠ�y��YQ��/���7܀%>q�y;h	�A�]��F��%.�lv��u��N����@G7���/و����n�nP�"��RT\������t;��.]�vM"�"3B�I�����2~  ���۽{�0����<��(���s,�����t:?H[N[H.j��׍S$�`�Ph&E�ӳI��
5�A����˯�t��X_�ՁFG�]YbB�~��[���K{���d�<r�7>�T�>~���MI��Ns�Bcҹy�llX:R���2��x �G�؆�4
�q�3e�67S~��l޼ς�9�4S\x�+WN�Ak�lqn`.�7���5 ]��V� .^�rŘ�����K�1�Q�?��N�R���[���Z�#ŐY�؀>� ��y����L��R*޸m۶;��/��/0|�_4��)d���n��)�!�1sc`����xa���em�%MA6�L��tu>�=���%~�� �`!k���6j�nRs�A~�iYG\,�կ�}Q��
M*�s�U$��_��W�2,'����jac��1E{|�F8?t�@> W���;z�bǨ��C`����ɡ��=��O>�TRm������X�i��[=l|>q�@φ���BK(p��qff�
�|_joK,W^�Iɵ�mN���md+d�f�y�{�B���el�֠rH<S=�2,�0�x��G�?h�>-�I^?mO�>�'~��(&q�q�@jx
�	O*��/���,���"�-��i����ӖY��tXh�Y
�|}�S��w��Q�?r�A����r)-$�p�� �����|�3;w���x�:�C���h
�}ۘ2!�5HU� Ǣ��>�'}��V�Ŧ��4�S�c9@"օb>�)�#C2���ӛ�UI ��B̡���l��]�N�bH>�GM�f����9�g��0���Ggb2&\�H��㬩�,�"h��yh{�k���߸���˼� �څl�d��zU߲�ME3�jd�~e�_��@�� KF�X�w��+3��Zg���YؕӚ�i����*�W�A���B�{��OAVM���[��#���K�D������?~饗�w�P�T1��1PM��}�=h�b<Ϗ�㧞z�^P�k�d��E��rU0�H�RS�L-�W��ՉS�%.S�^/�򐒦b<|d�Rg�g�>���bi��N�:�z���w&	6�Rk�<�� 1�ܡDͨ��گ��R-���5PC��r�K�P/�U2� �d𪖪�*�G2 ��!Hl����zL�Y11^��ƺE�}�v��9h{	�p�dsK��\���.�L��{���e�f�t@F͡2*�I^���E�ɩ���"66�j-IR��������O<�S�#8�9gO�V,󞑦��� $�D���ɨ�`��9�S4ń��?ss3r0d]��9M�ȸ]!����W^y%��~�%E3�#6z?��w��z�斒*�!�6q#�_�>ȥS�k�u��>����F�g�ķ�t�����kN'i���X��O���_M}(	�*L#�	v��;R���Ԋ��ol�YI�E��3S��m�_Kt{
%�����!>uT��s�b�EM�1NC��ZH�!@$i�J*M�"FԚ4�K�B�)�&�)yc�4]�����@��T�������j"olG�d���h���@0�	��o!'3[��I���/|h8_����;���z�bbG�%�m����: ���w�:���,boB�'&��p;L���}��Ǯ��s��V��{�
�J���R���-<HO����q$� ��'����3+&S,\���N�_���X-��Yٓ��~��=�u�0�VF��4�ÃXKSVȺ�/���7�,�8�D/�G��35#r�K�D��B�����~T�U	�׆�t��b�n��˪���]P��K�w*�҉V�C�6�a�޽����\p(��XwqE6��y?�e �I^����@ͬ���yM�3M"�4q�,������I��Ir�gF9�� ���$���e�����އ�Mhb&g.�.��0�1�Tp=p���w�y�E�����{�/4� �E�V*N�����E9��X��MU�x�h�˂$ ����+Y]^ޣH�h~v��Q.�������l���Ar7&���B�B#,���>}��9�IFf�/9ᆏ$r¢��'��$ߠJ@T��93��ZeD�Eq���P�8�h_��"��HC�Z���*#Z^�LL�9r	F0#x�Wм��k��!�W���H�0}\)4-����.��O�w��<�?�����㢋/xӛ�d�s����z���m$�E� ����xJ[�Ȅ�M
�̏[�����Rh�l&D�v��
q����©r�|���=q����I��&�ɼ(bi&7���X�.ҿ��^��}���V�����mKd�[�qc~��yf��m�Qj#����t���Ȃ�	U%���e˖��~��߼v�*�%�"��l�mR`�X>33'��W�?���b_�H>�#D~��1��io)	���0�}i�%�p��k�Ds-ʆ���rMJ��e�1J��-[��N4K�X����٘S��=�裏<��o��o`���G����2Q�z̨�J��ܢ����g]k_u��2Θ��=u�ر'�x�Z�֭[���MX>�W_}���iS:������,+�W^yE\A�n'7���E*=�2����?ޅ�X\��KF�sM*N&�.1K$�:oK�;ϴ*K��\J+
fUm9LgTs-K�)�zHM�&t��U�9�\$�=�\a �5 ��y�f��4�˶a�u�� �0�q�P�x�d�W��F��0�o�0����X��m���w�}ŶU�a9ѐ�%?��S?�я�;�<`nJYl�}���|��X�pm	���$��}�{�nd�i��&<�[�?�_�X��p�z��bM3i �)���~������o?���̛���쯴�q.�$R]N���mܸ�׃>��/�=�8"W�e�<o�ݨ2��D�Y�G�lt���J6,�xfCc��I�u����b'
LB��K~���a7��mXȐlc�^
��0����\�g�Ά��ќ8�*��fi�ukW�i#ü�t�<l�- ���<�9F�be^�,��(�DsL���h��(ZR텨�jŊI���fرc�˫NL"�[������vB!�i>$�>a� ��3���s�6h���l�C
���������wз����|�ͫV��(��}���vϭ�~��|'�]T��������G���o�V~�d�}|��o��6o�L�(��������������?�i9] �f����k�j�Nބv5v��br��:o*=h�^?E�Pkz񫛄��2?JH��5'�6M4I^���-�m1g��~��`�n3�)Zt]I�����GX����AC�5�z҂]ց7��VG���x��>�yÆY��X�MEP�	Cdl�� X����!%Y�ff�d��#������U
�D`��T9�T�-������\�u���C�� ����j��9B��RS^Y��	A<��V�/��{�]w�u��� y <��S�{���^x��@��x��"����4�Zs�+��SI4Ȋ���YĠ�i� ���u׷OΜ|��޷j�To~Ȉ�X�j=���=���O�c��'��:Z4VL-�.�5�j�O���Y��L*1����e�%��z5��v�S��R��SJm�p�c��"dYN�Ԇ_�;O>�$tLȧx#�	��s��_��_����/��s��x������
,"��m�q�T
���6������Sf�:Oͼ?r,v�{����-#y�;���ɟ>��r`�/���O}�����_�b]�ܓ*#fIJ}��g�����Y��o}+�
}ػ��/��?����C������|���>��O�˱G����_��o��� �{���B��9O+w��6�j��m�a�Q4TO�QS�;�i����%�p��r�.١������<b���	^A��ԜLV�zOT��*���ff��%��p��&̉�4-΀%F���,?
�O�A������߁W`��]wݛ��FR��ڠ�O��G�@�<d��K/��TՇ�oJ�t�K����5��(�W��W7�EEz�0�)C8L��Ca���~�M+V�Z#Ԑ�h��J:����F���c×��2+��ⷱ��ZK��1��Zc�O���pϽa�@vG��22����Ç�V�Z�a8X��+����Ӹa��D��^ݟ�5��sb��n��g�hҡ�Si((E�\�L��=-�OA�v /�fZ��{����3�v��h�i�JlĬ%���B�S�B#X�������~���f��M����������o��V�::fiT�g�rIh�F��δN�.א�~�fF%�XPH�%��-oy�c�=�v6m��z�E]x�d{��M��,:%�?��n��ۿ���ׯG�SSI_����Z�zbq��|���x�!���Y�g��H�g�hà���y�/Wע}��0 ��)%���Am�f����Wݯ����N��*�C�|g�n�@���L%�a��Z�?ٟ�kL3���"��]iS����IsWy�%��P�+U�&��#�WA#a@ d?��;��,���/��c�!�J�\}���O?���G�byKV��Ԩ�)��/7:|��{�8a����g���LT��BPgs�/��2�{�G���\z�L6o��m:AB����=�`bZ:�2� ��IRL��FU�r�ǘN#t[�7V%|����D�X�I�f���G�5�׻�����[���g~��C�<�}���[�ƺN:����|vn~rre:��7YI�x��j����]BX�ip�@���
��Zm���8S�+����bxmfbn'�R�oSҹ[�([�n�馛n��}���'w�n��� �{����؊���crӱ�f?�l8+�P�ַ�Rp�H�-6&G����nˤ�ܐ�gR�|�=Yhm����vI�:��޾m�'>�	�M�Ju�� ��c�- �#�<������,��1�G����A���3����o�� �׬a�e���fb|ji1�c� "���tn7��
T�=�n
�a�Is�`�5҈����{�u��[�͈�k�� �C��Y�b"ȴ���ic	���s�I�f�8����&��B�iQ��+8cwz�a�?q���C��eN��h`��U�"��N��=�܋�w��\w�� `�����I)�eS�[@?BJJr��Y�ٺ�\��MQݎ�X��L��P�������V��R�<��"�yp ��k�|���'sALG�P�{���&�&��&C����>��y`�Gߒ��z�[p��'�e�ڄ�b��B1�I����>�l��{�E:�!�����%�LM�ǐ���bS,\hG�ꗴ&�6����ť��5fH�
�pX�	,k��88��2u�2�2s
��.n�s�9��w��D|F��^X�m۶=��G K����~ݳg�{����.��VZ;�4IP�v,]¢ r�75�6R�����ՅZ/�w��fE*��Z���r�Oh��@�%`�.��?���~�~	��=�����7=rT]HT�J����trH)�I/��[��K sʻ����6L+�JеPV
�4�΂�XՀ��٬��j�̄(��m�z�2����,�Tc6��3Zi�L�̉|#[[���:�O��A��26�/|
<�oL.���Xp��De�i�;��G8ρlɌ!��B3�|� �3�<������8�/6o�L��˹0�����{�a20Kisɒ,K�:�əD,��6^����Av�D�����(.&rLl�)�1�센XXZ��>��sϿ����v�+Td��ɉ�U�fG���ƐVGM!Y��dʋ_�0"��c"$�τ��)�@(R�Q���i���ґv��������9<q�4�han�Պ�5�vn��9ȁ�sR7�j{�%��`u9;RC$:����K��2A�ls�嚤D�ڨ�mT��N� g��g
$_�"��J��o�@�^z9=���s��3�T�60o<������O�ӻw��ަ��<C��,A	h-����an6��$�si.qFГ���0��$�f���z.,��K#h�w��j	�c�����`q�������Z%ə�k�;��V2���Z
��.�p����r�TSzz��"��tE�j=C�(���#ցBK�s\�Ep��f2-�A
sf��їʨAS�
=�ͬ�|���zL��Мkެm=Z��z����P$��A�!���hҊG�q
�EN�]i�i��4r��J�3��s������o|������5k8E,�[j�0� -���e��'����+����������O3��Z���4D/�U%Z�,W��>8Pd��-8ٰ�Xb��{�5��pX��\h�p��A�8z�(S��u�/p|Rb~SM-io��h��7� H�}-�`�iͶlM']�)���jq��#G�����i;�� �KzV�e7P��p�"㊍72���<Ǐ�d�q%tF�:`�*��e��_����[>��OBG!
�
-f!�{#������ns\a.�ͅ�2�~�㊢�W���-lԈ�j"'��AH�	7m�T�Z�� @wpXW�1с�5fk�}a:M��؂F��v��
=��>�{�6>U�PH�/�G���p��&j0kx�y"4p'U�)�DgD%�3�5s�ƕKc��%c��f�{]�J��h��D/���soDgvkm�e�l�l���1΄MM.����(��MFl���>���]�Ъ�Q2�@��Ⓒ>k9�:��x?\t�{ Gdj�\цzPHzy�5nٚG�j��us<���lѨ}i� ��!�ބ�v�Z(�X�vP�����HU���}��U�r��L:�2e3eGP��<�L�!XK��Ƀ*�K>�E�J�M���}���9���r%GRv��?Jd��n�`���Z��r��~��D�я~�կ~��������=��*-�g2Q��������Q���'O���W������>	�z���`�����\5�2U�;(�`D�:�bq)�����_�M4���*M[�s;w��*eZ�������;���!��aԽ�w�L���9�%7A'OǽO���3�SĤ�;�e�� ��Ō�k�l�U��%�$2g�4�ݺ����ծȌm����$&Ǫ/Bc�E��A]�}�
�Hd=�Tްy�F~�a�\�n10��a��#�
OQ�rO�.��B+bש�و-��=�f�J/m�;�C�(�E���5�Y5��+���x�/:���7��<�{�(��eٷ���_�����|��(j�:��!�
A k������tCQ)f�K�QB,��ɔN�)��0�\���֭3�7I�����v�[����t���c蒭��L�2�	r�Kay� �z�	nVb	�a����ʞ={�=�\�©I�NJ3e� qv��c[�� M-��`b��O=S�dn^ǝ�J�*4!)=�C=�lX�Xtlzz��W`3&	�s�=w��᫮�ʎn����ђ����0ifq���V�칌y�f�Rָ�2[��������ۆ&\{
�6��Y��q۪~�x�Tk�1���d��V@��)
��'���G��z�ނ�V� ���oΛAjl���i�����솁�;reN���\�2���
g��\���'�2�������a��
#�4}�'���k΀t-�0�4<R�{�gp��^���|Y#�9Ù/���y͋��Yǎc���h�,���9&1S�H���tS�*��>���=�w�^4��l��I��.��}�e����ܜ��1QV�����霰PA�ǿ��G��̞bTP^ޕ�XAj~��ǹ[n��m۶�8��Ue�6۹s��?�q���K����{���.��÷�;V.��Z�l���JC�h)�H��l�&+]��0A!6�e�4&f,rfe���s��@8H��3��4��7�ꪵ�4��gb�رc�e�]v�ȑ|�Dh������mx�ᇟy�+�������,�\� ��as�9��K��Y��j���&:E8��;ԍ��Ѐ� (ƀ<P��U-��K*v�Q��M�1-�l��1F�eL���сl6q}��6i��H+��v�Dn2b��8�6$ý�~��ۿ���0��~���Ş�+�8k_ڳ��t<�x�{�||�T�i�J��T�Q�k�q�,|c��#(���в<��9yat��>�i�Z*$���`����0�H�sÆ���W_�����0W+0��1�Qӑ�c$Ǿ�>~�xa���u=-�Ƭ���%���Qh]���ϞI��smb�� A�PHD�ƍY�����ԏ>��]w݅;/���|�~�r��"��n���v�ͤNU�W�߿��?�!�����=o{�ۚ������y]��@)���1�r�U�rgۍzFe��Ӹ�3��q�i���;Ez�Z�Ba�\>6E?��>���ɱ�����˿��?��?ݴi��
�lh�U��c��m�� �_k���H�Unp֧��)9�j�l��qh30�?�o�Lo��F4�0�&l��lߘ��}]=�vy4�t�oƥ�(�Ʈ�$���Χ�ĽM�E
V� j�gف�p)8e��-��و�mm�.�����%�&�QQ.6_�#Y���DJ~)��$��z�rC��_{ʿ,S�#Ƭ^Π\Z��a��&�5/�r�pf�nݠ�h#�[����s�9� 1H�7������'�F�Hqc�Eq֕�<$�T!o�4}��A��'𬕔��xipU�����z:W�,�����$Q:�_ꩧ�8�I�:����<��v8K�]w"Z�S��Z\��`��Z�����ޥ��M7݄9��O~B37�8�ѣ�;vl����tE*jX�Bk�9 ���_��{��	�,p׮��<�V�a9$=�Nת�?�0�F��W$�rA�+%��*�������������M��XZL��0�L��� [�l�O�'&D�����k_��_���5�3�*sip�T3�����N���EY�A⢜�d�#�:��@#�Ժl�f�١\"x����I��ʅ好���7��~��^�U��B}�R6b�6;=%tW��W^i�����l�,[��/\Y�A�@������y;��(P����RԂ�Q���z�1hn�Q�~��@��cB��j�A��m�6�7fK����'�5��5�X��4�����3 ����˸��џ�cg����_J@�ȑ�'N���:�_�̄����vK!G���}�/�C"剱q|ƶ��ɷ`o3͉>:��f�*�	��S2��'�s9����5��dR�w�ݻ�ـ����^~�e0D���.��}�{~:��s�a��'UW�C���>��ϣ}���@|�O}��o�nJ�R��	�gp)���C�Y������=�q��A	��kG�yrʴ�K~�����W���B{@�R ����%�
�҅^��O|:~}��'�����]�v�����/|᳟�,������ַ�%E�����Č���[��[`+��o��If��n�t�m�ݶu�V�
����	=�~��^�z���������_�o��˂U��h��C�����Im�Q7'*陲<��9$���V�.���p�j����Jϑj��n.��d�t��Kk�
(�'|�!fM}��*K�!%E��@M�΋&���I<
�F���x��G�eQ�p���[� �I[�V�����j!~��}��Z�1�����7�iϞ=���f�с�s���9�s]�=1�@�G������\���ꅶ�~%∭ƾ����Z���ɘ�\�� �f)�4��M}�3NU�CJ��x�Z�7RI�ԫ����W��1��Z�z˖�C�G�vO[$<��� Ge)wgr2�o��������+&����z�;	�߫�1�{���5׼�[�׋� D�j�_�`�L�S*��6m��?�#`.�JM����c�� Wj�$JL���]~ť����S8�ف�<8J��%Z���9В1%}-��/�"c�N.���Ǐ^x�������y�����M�x:�h�j�Cs6���ox��߻f�:�Z_3�qÕW^	6��;u�?�K��;�Ʌg_zi�5ڤ������~��S'O[r
=�`x�L�!;߻w7V��v������ϫV�@��\<�M\B�e�sF�y\���3�])Z�>J�(�2����F���a�Wy�*�lvF�gD�Q0��م���#cɟ�l#���\���|�V"��2"{0=�#�R-R�-B��{(;86Yd���ы���pY�%�� r��Q�����x��E��8��:�YckJ�ӳ4���Ky�����h�����B*�\������� �c�*D��1�?���ʨ�pIe�F[϶@�����3I��(��?Mo��h��Ȑ�$�oR��5��	d����53I[��&wQ�b�����ZC>��`��͞9�8�~/�x���t�b������Z/I|7���jcc�L/��5�R�D�l���o�k�+��L�]����Ħb� 0�Ѳ�����[2���W<�d6�
��_.��4C%��d�ߒ��~����塟� �LuDʗW �ng���|������3��{J���k�F�!�[ O��~r�.������x����٥rU��i�������i�$�RO,jh29����w�{����L��zW�����5c���3���t*��Յι%I>p�:���U{`������bO��W�,9wZ6
�"Fv�o���,����3�/�&��?�4N�� �;������@�@�ڥ��=ݔ�Y.�#ˆdm��b��ظ?��9c��a�H��^�S^2w�_s��T4'�6f5��-%U.+��s��R�X�& x���2$ˢ[�� �֭i�-]I���.��=L�z�����r\���A-�x�*�ŧ|�)*m��ni�����|�	u���GŬ��c����/�v���|��#��`W��,��n�Ư���ǵ��N��9~�8��F��_0w�+&��D�k�f� ���G����(��A4�ǩv�h�	Y�Bh�i���� ���� jMȣY02Wx �s��TJ=������� b3fb���0��e��� k)vv'�Ьk���B��s�Bpв
�+-�^E��B���S5;��mO�t.n�"�h\׃a+ay��o@,r���3/h��dߦ�w�6[��[<[�(Ժ߿�>��1ڬA���w��/}�K 8���錨�Z�pZ�|�N������$_�h��7,7ݭoZ���fpin����=��I,���y�� ֣G�ɮ�[�n�� �7n�TW0����vQ�F)Ʈ;�5��ۓ�#7��K�H�$�<o�CH�N�h�Қ�:O�;�o��6+Ղ�yaG����}=�C΍��^t��@�Ql߂�s���E$�)��=��e>ӿ�Ma����D�aX��Ѓ�,���h���6��B ���gx�lpCW\���vj�����+�C�jy��P�VD⹎���7�i�2MV�I|���0ʸ8y��h����O�
�Vd��>�]&��yX�f���؉9�3ؙLe^�j+�Xh��Z�c!�A2��Ӝp(C.h���[R%n��+S�]?X�,���_-�k����-L�/�Wg��dtclVy�S��9Ab5DlL����߁L��5�#W���_�$_�9�Wt�L��3�',g����2�fN=�5ߏB
-!e�av&I��`�C2$yv8�*�]R�]�v!qs��6�'VUeI(�oM�J���oO]�rFkD��)�%�N��A|�F��"��B��B�^1��6)�Lj��5�ϝ̈F���֤�D�p	F�&�!�ZTXe��������)I�p�wJwxJГ�x����<,��^�)�e�7����)�X;z����fS<O��M�zKM֫e�$�J'=v�kJ���J��e�vdκd�o6?K��rb�)e�X���I��D�b�\��I������6s3Z� ��H+�T�RG�;痼��<�5�L~��bcm�Q�mr�?�$��9��b����<���ZPjnp�"��\�f�N��9���/�N|��ג�<�����-����m�5{��a���S5'��[�#G�|���=z��?��?���Z���:Z���u�Syd���o]�ٛH����#>����Sj�-ͷ0�CI�	Ɯl޼y߾}� �AY���Jgb�5)�q�n����õz�A��h0��Lm�9��Ro���aSL�a"*�O4�s��I �N�
���X��<]k���g�ё�f	I 1��`&#���x 3����ھ�T^Ru_Uޫr9���Kn��!N%�c'���1` a23c�I�HB��|N���o��Ww�s �k�p���k��������?PR�G
�Z(J8 ���.���v��L�~����C��O���2-|N�"��-�+�%q�c=
��_yKg�Y�;ƀ��m2&�����$S��b�f��mU"�Ji
W?=�S˃B�\��]� ����m�p��˄9�v�gͺ�M`6AX��
5A3���p_D>�^��qaңB�}��!�|ء�!V!��Щ��E��PvE<!�&�[o�t�z�ǁ�b���{�^�O�5����R0�U�Zە6x�m����u�����őm'�	�,��q>>�Olݺu˖-�m�h5�c��i�҆����ϲ#��7sM(��Lǀ�5+������[�L��Ā[�5�Ł�v��M��D[_;��M	2t���gw�W�5�.��)���rC+��u5r��>m8������)���w���<8�jhݹ�ԨjU�m=7bjϥ+WX�;���N�x�Ttm��_���IE�inf�u,��)����u�3]B�X|Eb	Ѯ����ߦI�U�J�bLJӁ��\�4��Lj]���W�����A�k58��S�3tM��#��)����I�g������SC���y�Ơ��V&W�-��0��m�_lD=��Oڧ�4�	��ΠX��b6��Q��W�3�����\�[���W�;�tN���'Aq�����p�J��Yo�`��[����?�Np�ڢ�q����;k��u�|�0(��"�Z.S�z�^:��&{��W�z�?�0g+���zx3����M�X<�yF?�Hu�s��]Yɩ#q�"�b��r���J ݐ+/�Qy,���:U�x``�x=5�d���O�>X�� 1֥����g����H`r�=��l��gP�i�7�j��[�-钲>���iB;G̢�-�B8;�M#xV���M�����Ư���K��!���!��Fo��U�����(�"��[���[����ͱ娒�w�7ՌN�Yz�hB>)�� �=<��o����Ap$����|���&�8�e@lKeZw�R���@��b�OM�V]�$
iP],�9�/>i�6�»�[u0�}"�Oi�h��薇if����ꙧ^��m�=D��+���*lg.܆� 	���|'�h�̬"Aw�J�(	������Lc��u��]|��b@6�Cr=�'fd�cZn8LyGa�}�C�i���cQ
��G
�%�>r[�ش��6%ڥ8H�h�bY��H�B j���T�.E�2f�Z�3u�37=UV����ѯU{�,YB.W�i�ML:��/j���U��<��#�?�<4J��N�e>eo�3�U+לx���Q����N(m��T@9WP���xwbnZ���(�h+O|��8i���	��-��&��p�(�f���%�,�j�Q˕�^}:�B֜��Vhu�lGAV�u#����/���ʕ+�C��g�\FoHt��߷P'�ZID��%zX���O�*��5���8x�o�	��O��O%<���|Һ/'��x\��?"�������=��e뢋.*����g!
����8n||�|4)���G�5��灉�D����L1�Y���nb����g�*�eREK�ꎂL�l�?�e����H�m�ّr��\nB�EQ�h:g}�����ېV�'ھ q����"�@�b�*��+Vh#��,�8��֯_�`���nF"�x�d�zv+���zEA^��5�r�g>y��i���̻y��D8��'�����!�T}����G&;�$��N
S��TQ���##�+t���n�7��a�''���Dm�[�-���+�<��s@�N<nÆT�3��'��u�m_���*��3K��3��}s���r+
��X�%�UX9Rc��q�3��������l��3�^��FO�ߔ����՛��z=F�P/0�ԩ�0�����w��`%���������uU�x�;v��S���{���/.Z�o�>_z�<�v��k���R)� Sm-U�ħ��!eo��f�g�y��s��$��mU�DA���L��Ü>����;�n��p�-[��Z����/� ����*�H}�$�j1#��4t@�`!��j�Ƚ�����Y�bg%l*ʐr����#����vE� �!q.��j'o+3ty��3(�ֳ;7�|��^�����K0l���w�¢a��L� �p�	��c=�sH��3_��dS?�����f������C�;�f��[U����1�Ok:�ެ-[߲�dM��^"�bI>�}Eܳ��E)v�fuzeH>��(I'?���V���ϥ��[d.q�M�?���£>��jO��n�ם�5�}���;w��+��'?}��'�;jzf��������_C���K�G�C�T�ԌY�V�,ȢƧS�)I���Y<u���^!vӳ�9UTޫ�AU�<y��P�f�I@^+]|W���ؚ�ӱؔ=ad�bs��$����"��Y:� ���p��?�'?�	V5��ly�g�y�i�N?�t�k�t��nֱ���z��k)qY��/J�W"W��yܶm����I�JG2%�}"�3�qui���8X ###�n|r�G�c�ҹб%�2�
5K%+�2�K�ϫ�E�}�3�
�,�y�]?�Ī6C�<�1�ǝ��^���Ŗ���{�X��L�~^62?8��@B��Ľ?�B묬���C����"��׬Ys��W�s@6YU՗
���2�j�y�=n�Q�|�>�ɤ�b�B��´6nm�e�2�B�����T#I8��YcL*R��d���!s���!��ά��?2*U�V�1���r�c�dӔ[�;�)����������K/A�r�!lDc:�Vk�*�j9!��8�DXQ/Ķ�ļ�{��n-[����= �A�7�G����C����Oy@v�]%�bM>�x}&�	U�Qy��3�����}��G%o%��>��3E���]���W�޽kى�@���FX����LF4��i�>ꨣ����o��C�gQ��-��R��N���O�V[�5K�,���K/��b�����zR�n�r))���J�����rj�v��L��r�M so�ҵng�U�AF҂�~G�y��	X�4�s/羒�*���q+���1��c�����Z{W0h� (e��U����Uf�I%C<��ڵk?��c���n�;: �@��mc!o$"�ݜ;>�-��|f�͢�	��6~��[���c�6�;�8(�<��)��Sf�H<|�e���.W�Ԟ���u\�}@�*}���r|�!��ɞR�RCM��fM#���3��щ��AG{k=`^�-O���}�P�q����&|�����}Q�q�B(s�7��j%3߷&S%����<+��'N1��a�"��K�C]�E��X���w$b
qkYz_e��/�m}}t
�H*,0���Dx���^���$�A>Ja��m��Q�Y�S�Q���zKW�ʀ�)���SU�*���)�L�þt�RB����*�u�}�7�qFr�i�ć/�ϔ���j���e��p����x��4�*��Vj4�Y�3�z�g[�+])��l��\�4$~CA�Pq�C'�vj����Y�$�����;�l�I8,&I�u�95��Ϟ={"9�X�x�%�\�I��h Ois7���A�P~�͌R0>�1�	ì������������O��b�
��C$��J�Ϊ��h��v�֭S�tzt0��7+8.�^�����ۊ����"_G��g���Qhe�`Oޝ�Gg����MZ?�kݳ�N{%�w2 �xҞn�{�;�Fp/z���ӆ��-�r<�%�TMV(�j�Sp��WI��˭q4�y�Mu��^�ׄ'=X��fN��}�!��6�S,� �fB��;wb����ꫯ��.[�lbb��zjJ(t�7�aU��Q��t>!Gf�s_+5t�P��418��g2}*L��b�/&�U��64w�`���3L57S��e�OQ���ו�I+CM��wZ�Bm��c	}o|�ySa�u�(���~���C���JEkc�mP*гB��6Ĝ��C0�čY[A�S'�|�		Ũ�U$f�����{�nU�~�C�y�P!i��laG�����%"=�j�1B3�xz�a�������\S����_�4�#�.Dm5"���$��Z���^��o�
o܊�9O����"4���PgԵE�� %�����Ҕ��]��@�M��N~��!P�5��4�8p��$�a �����~n��mܸ�0Z��y1v�Szz���o�z{��G	��	=��C�����Hr��n��
��c1٤�<�į7��6���<k��r�_��]���S���U_j�l�ܟ��R�7��"=���Ϳ��/���o�ɟ��)�����W��{߽��9�o���X�Y&)R#��cdzz��]٢�y ��I��X�p�_�!������Ie-Z�t�-���͛7SlC=���������|dժUt9��b�����7|�r�� Z��ԅ���/4�!L��ŉP��������f��>T�zc��5}�$tSp=۠,��"��m�r�!��547���nd/�o�t �������âݜ�N�ß����_a�
�akI�h��@���"dcR�]v>��o~ü
i�����Ŗ�Z��6�0�V�X�y�o�!^O�N�Լ�% ��V�@(O��`֪�X����"gj�\�n��|�4~��2�Rh;�2S�WW��g���AyaL�������� ����}��������i�֭��.��?���}xx�����~���<���j��������K/�Ep���_�<%�w����G�/~��7�����}hr�J��)�e��J���x��X�=���>�t�r</�����d�RO��O<묳XO�%�	+]tњ��u��9�3�)(�ڶ�I�6��'��o�>\ �����_u�U�q�m�f��3�Ԑv�>��o�[����A�<:��X�Oo	Z��n��ң�>J�ŕt�� �FO�������O^q�h
ψ��@��7���g������ig#s��l��Pr�R���s��I�	�y��%�#�˗/�H ��Zc}�x�'�J�cy�)w��TνO�zop�R����� o�)�d'�] �2^��veHNC���7���AŇ����7~�(2ʯ;o�N`�������z6�pq�ǯ�DR��^��jH3VdUWgYXd5rSTsq��%��EUH6C宅	��J���F����`�7��J�'6���鱑Ѯ�J�鱦B���E�;�Ѫ���7��v�t�(+j���~ۈ�\�j錳�L0���uQJB`��Vm�0դ��@��g��L�qu��K�7zz�֯_��3ό���<�N������_�������<3㤴�p��퍭��4� �6*�ݽ��	P�������_� ��g���W������z�����o���������f���BPN`�����Pe��"�җ�������k׮3�<sl|��[oŇ_��O?�ԫ���%�����R_{�xj �䤣��� ���G��ڵkAf1'��vǮ]{.��s�=7M�������[�� ڀb�����2!�t��n�ڮnǬ'���$�h73�7��sn$.gJi�w�U:U`!�4�s���m��!�
���YP��ǦH�^�������7�x�N@�{쉭[�b�%��4����;�m��'�,�h!����ޑ�	ܿ^ϙk>m3��SO=��X�ry"�n�J�e���^���E���Qp�N�l�H��q ��(L���a:Ϩ����zkzzwy��$p�9��?��O~�����S�F)GC�@�����]���p
:Ĳ��J}��@P�SxU�g�U�H����]�O%�� e�<͢.R���g�իV�Z�\3ˍm���o��VC�+��f��Nn���5�Ty�3"�$�	��&qd�>$����m�<�1�z���ʕ+��@P��Y� ��T���{���{�^{��y��Q�-��VE���炣oiGBA40��͒ҥaK�SmQ��&Ay�6q:�P���g��τcj�/ŏ��A+
��ϥU�*��2�0Z�	-y�K�3ou��z�R�>/�C�����O3.�|v��� qag��R�K������ݺu�6�!����g?�-6~~�����q%~2::�@���.�P#L/,����=����w���}��އPK -�pp_r�%�u޶mP�S����_��M�x��(4�Ï8z�� ��=�܃�h
"��&�:�nŘ�jP�sO�̆z��K�~�-OG]w(��8��X�lw���j��\s�5�^z)�,7�|3dϧ?��#�<?aI����_������_�j���/�p���tg�z����O��Úƍ�O?����l#l�A���5��������A�:��b1��{�H}���5����g�P��'>}�mjx5���T�Ž�Ʌk��b*i<�EA�����Kw"_$�m�`݀*�"�hI�=���p1����9I/��w����v��͉�����O�FG\ջ��˗]z��n��Fw�=>#�fyQ��R~.�`j��T�!<$1���ݞ��\�Y��� ������e�����dTh8�1c��
hzmr�Q[X�a�8^R�ڬ[���F����)چI[SL����|�{?*�C�t��O5y^d����[��EN�̍�Y� Zᨣ�Zq�d�z�XAM�ۏw!4s�1P���b�/���o�$nӦM�mX�}�f���롇������^p�at"�JQ�����������Yg��Al��/��7��m�` k�c���v�mW_}55���I<0���_��'s����SDQ���	p	��g�gt�;�î��*����P�u��Y��REWQ��4x8L+-;�aq�r`�o2�{{����n���7߄����%���'@������p�W��x�L̥^3��EAɁ�7�x#^�KAN�L�6�DCBTw)��Zu����K��c�¥si�3,�$��M.���QqY�"����>�� Qv����~�\�Jmff�O<q�1�6o��J+:�7�<�ȯ~�+��@�����ܿq\&��|J/u)	�&�I��S/����4��2���K�_�/�Cms��m����ٕ�Q�7��E��y�é����_����'������k\Fp�}��]Þ�$�Yp�9� C��0�`@t`�%T"3Y�ËSV��EB�)b��ܖ���a�Ӥr15�e��fh c�b���2�M���C����t�_�Bא�T����bmA?	9uI�MS�	�Cn�m��`�����B&�I1�e�8}`y�� ,��Ҋ=	=�3rp�����6�c>X�s>��@p[|�J��/���� 8�L7h�%1�K�(��j����i'�6��F�n����~��W\�,��Z�c�!yP!\*T_ݑ�%h�#��!��Ǆ-`���$�*�T�مB��UMa�7�HðHt���0Dڃ>H?��x뭷�˿���˿��}�C�1B�?����P�|�+�뮻���o�[t��믇8ь4Z G<�U�p]�����A���ևJ2�m�+z��w)�:��F	�9餓��o��Ӵ��CA��� �9��r���z�G�t=�e
���Y7��d\���7�ǌ:��,�]��6��Ϻ���C��p�u�n�y��n�>�ęb6ӊ�-'����6���+�ƹ���T������<uZ���Ă�ڇ/������y������@�V#+G	�d2r��[|#�sI�(�Դ�SY��J�س�����N3Mx*�Ϻ-���cq51�]�e���Y�D��Y���d�<�9ta��ee�=d�a��(C/�>�?�g�N�ML�a8�iy,� �4��t#�I�Gn�#�»��, ���[�{�Rq���n[�Io�d��/���411u�M7b��3���: ���Ɩ-[xR��S|iPx�&�ey����6,XZ��/|��eX~�ر����4�PH6�����<2u��{��M��ȡ�D[�e��2�wtM۸q#��O�S�^�4T�na�:�B??t	}�M �D^h ��~<,��_�5+V��4�+��[!��x˚����d�h��E���J�m7~�J���
��ry�i]ln�r�ҋ[�`О~�Yp����->��㬉��r�Ú�k#���{��Ǫ�R�՚��@]_#d?Θ�3ƸG(R�2������a&��]�����y'/������|;�?�fV	�6�S��+@0:6�EI���J������*���n��t��/]���_m#��aa	K!��}<1�5�le����AH���;�g�J��%��\ϩ/N<=�5��-�G�&�v��'�)).oٶ����Ӗ��,��*����U%>n8*�+�24R�
t��� 	0h� �拌^�0�6�w�W?��n��Wh������~���^?�1�O�2���1��l��g��}�Ǥ�~t"� �{��^�����Y�}� �� a���hspp0�Ы7
�Fe����4�:Mte�]�x1h�<�g^C鄗��p��C�6j�z�J�B���ԊT�)�h?�L�>f�]��?�!�F>"�����9�)m̈́�fbJ��gbJ|�pz�QB��7�y��'��� �M/]�tŊUts�3m:��f��Tw�ܻ��Лfͨ�R�e>c_��� +���(�Ǿ��L��Z1̌:rL�:7+��B=�K�O��ě�T�{�l�]v�7XZN��~m�B�|EU�U��,�n;�o:9�lp��t�Փ��&F��EP���I�1��q�Q5�������	�J�f#�yjԭ�(u>F��<>��6]�}&^�	��5(�Jk�� �GHӆ�*�#��X-�5ı�.Jn������j��i딴�����"�Ѕ����
"�i��i�v����s������bz4}�
��Κdx�@�ZіI�]��"��Fa�'�8w��V�I���_�� �k�����N+����Z}�E��@�w��'T��\TcFhu�E^v�e,�6Yc�555�.3 Δ�� 3�ߍO��t�"�]A�Ng��2�gd䶯H�~q�E�5 ���g$�"I���٠�-q�)�D%�3�����^��j��5N�ˋksW<.�#�/!.��%N,ff���VJ�s$f�г
��@�MA������Jm�R�"��AP�M�+sͨ�7gVɜ�O�6�#���澢���)�{V]����N�l�V��wO�3;<<eH�m���M�n^���4>�H�U`�m`ik�2}�W�#�l`�aW0,H���([�(O�0�;w�X�]5���j�,��v/�쩕��k1RC�����̶Ƈ�a�:���g���*�e�&S���Α*Z���3nIU�}ds���-�~mиnr.�������Mg��\���q0��b��*`U��}w��yTұ�oE���K���o�����������.�~�v#�N���[��={��{6m*�[�]�#��Gǌ��0�BYw %S&Y�ݍ�����@y m�v@Q�nh_ː�o*(������/b���O���Cڢ���H?1��0���(j^C���'��2�JIC��Q���T}����b�!�៦���
��Y��)+q܈��2����*��h�S�}E�6��3	�_�j�I'�4==i�
5T=1��4|̈́��>��SBo{��,�[�g�	�)b8D��b���?q�B�M�Ⱦ�=D�wT�i��6d���m_!����m�������Α��~�@B"	�)�r[��\<=]_Г�|+{mxǓ�O{h���2LNE�*HV�E��b����4��˳k�GQ�<����ݪ���ٞ�V1����-�L�V�C��卨���[��L''��9S�˛5�3E=��e�ٽz��⬐�"�7�[xRh-��@����}�C���4�_���m�Z�>B��S���=�����l����뤬��w���~��M��Z�b>�'��U�L�xd[Y�z���nݺC=]:p� �y�57?��;��h����$�4ה��k�Ư �� F{`�`��5=�NՖ/_>88�>C��C�aP����n۶m��j��|%@��i�! �AZ���ȩݓ���A ��2I��c�X�0�7�Y��Gj4࿬˞��.:�O��׾}��^Bj��-x_�M���׮Xc%u�l���S�ԇ�o&��1���t�q֌�d�Ǎt*��kL�;�e�%�'vc"�C�����ا@p�FQ�4׍)뻧Jr#_�<�F�'<��셷�����>�(j��ʌv'b��Yhq����~��0�,� ���P�
1��M۫�UW�U~������-��tWF\`ն������޺�Ƒ����8��;���3�&��N�ʜMܹv��Pb�����4���"W/M�H�Z@x`�S��p���lӧ������څ3+�x�b K4��	��<k�~,�?Cύ6�_:����2q����c&�U��$STr��m�T�i'���1��!��<qꩧBJ$)@�t	���K�.uZs�
*�������g�u����0Exב����<�����.���|�{�Ûk����SN߿?�~������.��'?�I�	�`y7�t��ꪏ"��9���k��IxfZޔ��FD�~�a3_� �{��W���?��zHU@����\�k׮'�|�?���y�f��@J=��3����\v�eg�q�ڵk?���q�����S	 *1[���֤`薗�� LӮr�`�1�����g�$+xXZ��0pٌ��DЖ��^t�ypp@MIL���C��6��������w\�#�4Y��hj��N|?e�!���c�s~Ŭ�W)�*bv��\��oK�;|�W�y��"C�D�y�\/qg/� �E�����i}����vW�&��^3=����f`΢�bKQ#.�(�s.\�z��	}-�qU �LJ4��R.H�J}�$����.k���&=y�W���J�$���K�kMK.��7@O�L(�1xRO|�׌>�$j�3�u�S��5L��^��'M;{���^qk�)�#*��#��y��n݊� ��?�<Q�����n�x��/|aݺ� �޾n`%� ��U\u�UP����30��L����n�P�]wݚ5k���>�,��W_֣��<�����> �rr2��[�ɋ.���E�`Р��<�Xa�C�+W�ķ��V�[�g��׷�ܹ��K.a;�)'.V8e4ę���	B�Ԣj|�G`�7����2�e˖����݅G۸q#���u��C9�䷿��#�<r�QG���4����=�>�cb4�8�0kt��.x�խO?����>�����(���&&�y���Q��={v�w߽�w�(.	������W^�Jt����1����5h*]]UY �"�����Z���p�d��}�cx�)�y䑏=��
~r�%�y�H�e�|���}�c�i�Uʰ��R�Z?�K�����u�ݱ���TiJHVJ�fx����tJ�i��ҽYFΛb?������k.�5��uK�T���w�׹�#�3T�����y��r�!C�2�]Zz,T\�6IQz�V�$Y=����I��%���7Δz�.���0��P�\�-�!h��#�A�`�3������ȃx�#)F�s��Y\���'$��T�(�%��ZB0oI*A��񀿫W�.�x��֑$�{F�l]����O#�w���{��}��o��������@�+��rӦM P�5���Z��o���o{���q���g��x饗�q0��_@�I���Y j��?��?��oݺ͂u�C`1um7Y�+�W�Wh��o~���F��÷x�A<�����v��CPQa"��͵�r]3��N�;�3x@!>y�W �b��P i�A�:��-Y�d��>�h����>���8�4t9ǥJ/����� ���R<��(�`܂'(۶m��#4��Fg��΃G?�����&|��������![��PXDkE�8���yj�Ɲ��4����������	���'�x�+�@O�ϝ�8ʲ__���R�yI�HG�^���R���A�|Y����heZ����%YQWQ��y�J�Ҭ��ޙ'��!��^�C�e|'J�'�;%ƥC*�F%�m�a��ݻ�}c��y}dղ���X�}������"����L*~®�4s<�+�d6sKLwu7��Ta�����]�`.f/Z]1Պ������=�4�<v��jR�C=��-$��ڞ9
Eu����g�����b@K�����Z2=]���.%���+I��x���*�ui<�����7cIڀkN;�4�ҹʔeб��p���r(��p5�A�N�2�Y�j���G}4voW��@��N:�	�9\�~=���kfK�P��7��޴�H��`�@4pL��Y�M�z�N�L�PGv���h������a�`Kt��+���Px��c�<8dL�WD,ĸ��,��Y�>$]m��g��'�R�E�+: ��s�I9q;���n�i������g��qS����mƳ��_�5.���[������/����{rvHS&P]�x�^����"GFg0Λ7o�~8>2��ɸ1��_~�W��uI�҃>iz��v��ё�O����ʕ�1�IR����� �T���x����_�E��s�9묳�� ��F���g?���w�}����{{�9�2H��g�f�Rm�.���!%˲*�gi瞢%�{!��x��lI7�n��{yU�'0)3(q�o�}E`8���C��C�y;Ԟ�̕O�a�n��h��W޿g�:Vv!�!]"1�Of��ON/s^z�x�9��,��5q��^����nw�QHy�\��X�n�R��N]�����8������7A����*�E�'|Z�D��a\~dm[©j[p|�p�kH�
����W�� �)`1�biV�"���s}��/��8�ZB�*�+3����;u�M���]�n~���nͰR�|��NN��i#,�:gt{�"��v>��?�=M��Hg���=����"�=>j_����$C��P���ȅwN`�M��W;��O�N��#�1�?�%��!������}6r�b��ٜ^"h�3�`B>:����9M$�b�v^%���Ш[!F�a�ڵ�sgBqe��|��������A� ����y�{8ȸ~`��B�X1׋�tƳ����X�[2�g ���	�d	�-#ejV�g�ꑑw�
�[�K�L�}\����2j�֗UR�4�1�䨞��ڶ�:8O��aѡ�v^3Ϊ����z[���f��%���Kw`�Keմ���n��ܶ7��7���d����7ނ��fђ%�Ӛӌ�[1S���v�}�3���@�u��G����oa��Ǽ��Ը�.f,�jy#ߝN$�c���t�����Z��R����TM�h(�,�J��'/�_YP][*ow"�z�`�A0v&�'l*B
kө�����dA�*dX�����h�X�:ɂ_h�ӦAO�*vN`��� e�~��E���^�nK��]A@�֪H?�b:����9�]��t�fL9�N�9�G|�eѷ����f�z@L�Q��8�<���p��Zf�N�J�&0�3��]�ݐ���CP�1y7]/(�)��2�'�2:�%K�}����F�W���
F��7�9.�VY9��:��#�ȘqW�N���g�q�d�a�p�?opp�6<���_MLL��-��'>�H=!̳r��8��-�)����a׮]�
g�}6�C^�ʄw�2��E.8;�{_��yC=��7��� ��x��|�kȲ)�"1��떉Z]�������&��ܧ�ܨ���m):ߦ+� �����z �6�)-��I��ϭ�*���w���K��ҥi��˭�_|�E�4s�a;N8�=Nng
��r�#F�,�f>%R��j;��M�W�~�@�^߻�)�TI$v���k$!���th6�U��yڞ?d����/n����V�m�����U���e<ء',�6α�F�Ny֒ʠ�m(*L�!��!E0f��_��͍I���h���F� @�����?���/C��v�l�
�@�?�`$k��Cj��"2D��=�د�k����;��'��]���f"��5!8� Yk�|?�խ���Y�=j�k�1G�����qm�n}`t�˥>�U,q��Om����<��3����n�iY�(^��Xy
�b�*5��CCC�K����q��ˈ��ظ�p�����+�����]��8�?=Aƀk��
�6�A 
�:�A�ѱt���-���pY2}]�ϓ���,(^�;��}z<�e�vh��(�G�+��<͂d�6�[��M���h�4k��f�+��ߎ=]�L=�����6�o{u
���]M��h��';O�L[��6l�hcΝn�k�{+{�Fъ�Ch�n4VsL� ��pW����L�q��U��H#u��ń�(�v��{���P⢾~��9�Lx�C�%[Uփ�ת��a̲4_2fz+���M|-����V�y˔����E#q8��>*���/�2.����?
�gec�?@aZU�E`�в�Q�KY*��_@G�� �][�脅�۠�%K�QF����Eweh⨒��ݥ�bz]�RQ����#�ش�s���a�W�XM��m�;��UG���u��~k��� �qi�!���z�
�X�"�U&(��0x�pǌ%��.#�4k+�[�V�n��u�R~��$�>�&�"$x"<"E�lU����4���&�h�u|�F�HȫH�oZ�_5�*�[c����&�ɜ�EHYT�2�RM]��yȓb"�(�Rv��D�7B��n�gy��6�c�q��E��C���C�S�,��6Ѿ���2čk ���(oĔ��^H���^ʪ2�~�Q:�����8>�fơ�ӊR�{�Nݥ�UL3�b��#�i2_E���=��W���Br����#M�8�X��b���5��וĺTA.I��C,Xaʤ�22��m΢"��EC&��e�;��VZ�t��GB3s�c!��}��ߍ�N@׋;��	-����y\�}�ͻ'i�%���.�WYf���E@bD�� РiF��������v	d�,�\�J�2��a�v�Ǌ{o�_�9i�.V���P���>L+�śMkE�P��5jԘ��)��]Z�9��"��w��񞪺vCɝi=�En�@:9�i���:�e�eI*���ض8t������7rM�>�h�S_*Io�p�͗<��{�&D��yQč��C��÷�(�ʊ/�?��Y�Nc����I�T|�L��T�J�@�$(2k�A.%(�\�p���h�1�'_�3m_�$�vR_���[��5�.Ԟk�	�UjE��$�0ȃ��Q�9B��c$�П�R��(�
XR*7y�z�G����fz:#q�M�,�S(ix��hK��%��k)-^^�G:�:�z��g��c�� #�Xߟ���m9쒝͖b����J��.{�x���Q�7u���7�����m��._2�]R3fd���]���	}�j7���צ��q5�]����Ff��>������}��M,����q�'Q,1l٤��Y���`�&Fg�G��O���]�>�e�]���Φ��K���9������bʿ��df[z����d���2����qݏ\�=��\�������Q�Ovj��C�ȖV ����U+]��&4����G�qg*6�� C��c�����K'��Ҕ��Gm�,�1�F#��ِl�j�O�̑�ԝ�C���++c�K�i�UN��H|1��W�W�*���Ǝ��5|����n�Mu��8Kˤe��O5E�<�^`�U��K5�ܟ��3U�ͦwDy!@����;�s$�T:e�������#�LA�0~Bګ6t�u�b����S�2A�X2>�~�|�&�O���fD�-�b+�.ȳ�q˱�ӧ��M�VD�S���B9��u���#�X�U�vA�B
0����d@KX6D��p�ma�⾾������wo��=�7��ٳ}�v T�d7�qF�駟޵�-��E�j�x��1(��a�-��i��3�=+���L�r�N_v;��#��� �|5%�.*!�G �Wᔴ@��5��'�t�Fb��5�>G�,z4W�.ҕ�wT�����O�F��h#mϮ{��U���U9Z�X�z�Rr���?t�R+��g���rϒ�]�)	�	�����x�!�H^�IRZ���8J5�02��sq`�2_�WP�t�!��ɡ�~�7��NF4�)�,[�Fbg�EjXgS:e�}=���+���A�P�O�زNh��O�Q��6S_����F9H�Ӓ����2$>'��M���_���fU��EIV���MDRzm�'m��i��+�4=1�o4��J�k~���'�y��a8�j������C�OlR���oۿ���[K��(�M�-���qp���vlܸq<�1�z0U��7�7g3NO@/N��'wN�Yj��1]����W�|M2:���19:2~�@}j$�W���-�D�gK5/�6y�+&!'��$����+C�o8 ~������g\4��Bs�){t4�r�(��Z����ۗE���ǨPf��C��� ~�;��L]�G M��0'�6�2%���6�"�>���#A��MK� �ف�/�[��.߈w�PE�Z�*�<:r�3����툹�Q]�� tDZ����Ca���� Q�A[��x������CQH���^�nS�F" �+��Nr���$��|�\�-�V�)����2j0�m��>c��2�%��N����]#��X��I����-ț��|�,�ʑ�$*����Z�V/f��$����6����e�p��-�zY�G�|gt+�_Ȳ[_$��uҠK��=Z��B��Ƌ@����Z���f�9_��]���,W�Tn1����u���8-ґ�a�k�d<�U˩E��+.\�4�����dt@��U���|��D�L��р��_)�]��c�{���b�U3��&�Αj{
3�Xn����VQ=��0Ak-���(�YnM�Sb[��&�*��͋� b<�*�b^x��n���jT��4r�7[����B�Ѻu�`�bՎ�RsT%A��0W&*�5G�?�#�� ���r�yT8>�`=�WiǠzL�WX\|mV�&U�q�]���-bvU�V�΋�T��_T�W؍��5Q�Y�B3q����5�;��hƇjHfz"�^��p�*�5���e;E�0_L�[?J���R'hz�P;	gJ9{�<L ���Ż�-jqS��������w��hn�v['��%�����:�����v�pf����r%��dV�Z�����ې.**�T:��ͷ��`��V-�����O�3�R�Ѥ�{٢��7�|����a9H������.�I���˱g��j_�+��|��Vd�0�ܥ-o���"���lj�g����޾t`A��i%R%L�R�E!��O�L=��?�lb[�,�@b��
�I��k��:>1�]t;�g�+�$L�6w���0�T�!2Ƒ���a�(�$q���{%Dm#��8��Ӵ��PeVB�
�����S6Jd�
�������g��-T��W[j.�Q%jd�\�	��NR�J+����B�,������$=�,w�����VcW��(�ҍ3b��У�D� ��ό�ïk��/sV�Q�%.+2�J'��Қ$c��QG ��ZQ�i�0N��%󗾜W��9�z�R�ƫS��g�=i�P(E\�+'"��-�.���2L�V
>]�(~G����g���"��{���mx6�<^x)w�%W����H�`���1�H������pC<�R�"�V]���n��%�=X��K�m#�af�o�a�npL ���F��!��7"l��w��i��V�\9>�ϑ/Y��/�|�����ū�85�d�9}~]�T��Q�C5؉�Q�5q��冽U��bjz�ͺTBR�T痁�<˻�6|�HNzr�q��Zw�mMR�|!4,v>Z��� ��L}��7�}�F}|��E`NQص����gv�RE���
pz��'�[�*�)��*���d4�^#�|�@vF�3H��j�a�#k�X3G���b��ZRI.�΍7R�A�@Q�,+�u� ��1�z�e��6�U�N�*ӌȉe{�_��/5�W�/�F������mk �iH!\�W!u0R�+�qC�^�dd���f����H]�&�<8��S�pI�>��]�?�^"�U�P��������fA:\�ym�u�?�VO��o3��<�~<��v�F�C�d~�������MG�֢(�^��,M&�M���ݨ�Y��7�'gl�3F|�z�l{=˗-[�wϰCv�WX��i��5珚�ZQ33S���M�ǩ�Yݝ�W�d5����LCn<�݉�7����V�+V�jEƕ�������!wFcc� -?n�G��*�P���?�"�T�b_SNG�k��+�g$5���slט0en-�#���iw�k&�RI���������*w�u&q~��GY%`���kY�g����\�>HL���!��k��v����7*7Ԝ��'S���.4r��K�5�7��b�2"n&tJ#^�͖-[����y�S�}��H�W,�+
 yGvIlǩ��'E�]�엠 �`|Y,���ۅ7
s���cL��A�k�����u/���z�!M\vg�J�Yǝs�)�@�F�qW�\IV���x��-Z}4Y��R�^����C���x/��֨�t�*���Źt80�:hF>%��(}�D�PS��55:)R[_�H�L�xȜ�� f�U�+K�U`�d)1�QT8�FR!��(�[t��6T��ͼ\�h��J�������fi�_���w��������3�`�J׼^�D�cldbjp� 6���
��̸�fʞj��N21�½�E=�i���Z���y���⒅]�F���/��(��f=����y��GT��U�r�6�G�K��l�ݯ9$/�3�5i�/�7y}��idd���C-_��v�-�?�x�
�~��B�d�`�A1'�	t{饗�x�M�6q.��Hi��h��h�BRZ��S_�O7'�
����w�}7��/��/����R~X�`���|��7
9�\�`��W^�y��i���'�3��p�x���;�{�9�Sv����[;�?�|VMdڼ�vI1��sϡ�^sG��J}�E>ӧD�tV����g�?8���A�1RB�0��S˱�5��3��cN��[ǳ<��ø��O^�beث���9����S4@Sv*�σW�tזb��_=�(�xw=��I�ڑu�u��d��ā۟Z�ٱ(���'����Nr�'ݡz�ӶmCh��ۃ���S`�u�P�q��N>)ņ�;X5��A>,�޵���/>������_[sH%�O�MXdw�g�Q1���K�l�J{���+��≉�����dw�ֻ��E3&���.H�h8.kA��HB�#�J@���PK�jW��>ypr�@^_C�? ��V�p�Ȟ�ᛜXڂ�k�QE�Zai'jb��u��:�S]��8P����cEu��k��<-L���@l�6(�`���"�t	^�4�����я~���O��+^������c�\r	5;�����D�	CL��]����r:RVPڃ#�g��مMW"�G�XJ�%(�3I%vic����ʲ ]�"8%R�1�����LҰ^��� 6�j<55�a㡻v���/~��_����$�?�#�Q�p��R�u�]'�t�QG��F c�/�=W�*.7!~�t�R�Y�_~��Ø���Y=݈�F穧��o�9�>EZ�3QPI���������S�V�Z��\365A���; ��η�����?���E�w�^,�c�=6�t�hp۶m-$n�.�w��NI�,Lz5=��@N�ݷ���CW-^�x�e�����m��G�M%��\uViStu;��)�>�^Ԏ�<�M��[���"�`�������&�xaޚ�����E��+kV�[�]!��>*RC��f`WΚ;"W�C�C��
"nL�-=p:��}�'Xį�N�n��Y鶝�H�ւ�y���[���Q���;e���k�J�}��gw��UH�����"Ʋ>0�o߾���x��O&��Eԙq�m"�q�\����$�̟����U��K�.�������U]m��;��m��J�g��E��������լQ���!��Z=�u��~����{��5&P�� ���uT!�>�$��d)\�p�B�C�]��$|VH{��f>�G×k���'��u����iӑX w�y���={�>�?Ͽ�,�����	ڿ��K����ſa�#٬�U ���Z�2�I+� \ħ,v�M��x �Zu5Z�X��峠c��.+4��L{�>����ͯ~���d!g~(�6�-t{�6y�G���z<>�D��aaj��~���]w݆4���0���DN3����z�UW]�H��&�3�<��d��e(`8Ѭ���5
�I�]"��������Ub�t8$����B���z�kd��B+�*�������CSI�3nȊ��U$tBa1��@:!�mAf�?;5�YC'�����!nMv�y�{��k��-����ڲ��#w��\� \�@��q�Ԗ�۵��oŢE�T��z�Qz�hHW%����$���Xlcq��m��
���'�8lxl��JW�H�$5i=��0邸�\X3=/,����6�2�*L`�egL��?��)6y-��Z8C��G.F�FR���9Z|E!���o�`ӟ�q����r�
rj�T�MXM��7� j��:�K�4�E�Jf�B���m28�0�b��Ġ�	F���g|t� ۼy3����
hFx1��QG��| �(<�3�<�HP6|�S=]]ݵ��?��+���	�K��q�&f�4�ܹ�[n��\pP��p�Mh���^|�E\�����:).^O�H�. ğ}��hD��pD��k�b�t�BR\8�U�.a��n}uxx�֭[���*�t �Q �fb��TOO��7߼gϮ/|����h��Dp�+1�JY�Kc����}Xq���*��F��ڵk�չ�%�		����qCk�� �k�@$��))y�����Q���r,]�����D��N__���t�T�C{V1N�x`�_�_!��{�xsb���늵�=U�^�J��ۯMWK�����ȇ�Fj�T)b:�N�\�:�֌K$���{r���g�킟hF�%,��ڶ��K\d��]�	�m/��mdN?7����mS��S�B�dnZ�o�	�g>��'F������؊̕��&�QamӲ�'�%K��LL`G���H�tB�#��c-֣���:$�J躘�]6��<Ib�G�x�;���Ǥp͚5
^Nh�YF�Ζ����:'�����g��6x�9
q�7�� ��F�
�y�ȫ��/�:�*GΫ&槟~��g�Ňo��&f��\�뮻�9� �%T�_����{15@v��-�[����S�����??��߿���@"�e߂�5. ��NBB��;v�{�R�������n�W\?����|uH0R�et� ����?��ӷo������^�_|����� ��k�z�{�[���GS���g>������ƃ��׿��'tP��y��^���/<��M@�ݻ���O�g�����n��rt���pX^�֭������oĘ����g�y�i�MNLXc_�����SNY�r%:��<��1��w��`r��������?����,HA���ׯ�������+N�T�ɞLj�p��) 1bh���Ժ�x�	VO^�b����g�������Y��C.+s�����j�+iֱk�w���Rp��S]9�\��7B���՞�׾�h�߹Ui~���ö��6�nk��ͬ�ڶ|HW� �9jF���vi>�ֱ�=�>N������%�վ�뮮����W�vM�3<����3io�;vp��kǒE����6c��w>��-��<��D���S���q�wU�bk#�7�=���}.%q�D�J�98�at�y����^�~��K-h�<�uP~R����/�&�Z��^�7���#��E#�t���@�#(�DG.�H#-S9NJ{�p5%eJh�;x;�CX�����z+��	'�p�w������'?	t�0nڴ	�������{��7�x@l%��S�w`ܠ�O>��-[��� @�����k���|���_�����`p������J<�m��v�'�ڏ����?~m�ƍ�_��]�v��^��:\V|6h��� @~�A��qǝp��>����V�ڼ�}��k��r��Ǟz��5�S�^$��W��馝��^{-O� X���裏����Ra+g��w�yx^P�s�=�f���]Õ7�t�p��_|��Qj��}6��[1n�v�����)㿉�`���e˖Q����[�=��y�4rWGB�2�R�x�w�n�}�WB�A��+�H_�(.F��z��!°CO��_�q=-�͘��˗ӘCd�ԃ�C0]���S��d7G�i}f%&�4-�[m��(o���U�s��b����vB3�+�2��L�N�����-ߔCm�mKw�7�0�2����3���!��-�6��Ag1j�|�1i�_��fޭ=�M�"��m۶m<�<)K'�����u�$�-����Xy?�-�|f\�
j*F\D�q����3������n�r�5������M�m8/���֩�e@��<b΋�u�A�߲v�q:��}P3�*�F!,fU�R�A�.�.a�$��礖4��}���9`D4H����~�S������.��|.brd� ���� ���y�-�lذ�K_�>��8p_�"%ܾ};n��� ���ȣM4��4O��k��&�L&Hu��?�ɉ�'p�|�g �������}�� ����sι袋 �xF�x�����-�J@0�DN!� t��	"����?e$�_}�U�9H :z������TX�x	:O|����~�;fww�<QӶ�3�T��A����Fo! ݲ�*y����������T H0;�!��Nҥ=��{0��9�0<�&�|߾}DpZ䡗����p�u�AB��'?����?͔��o�l
{�x��%`��JܰL���Mg�������2��f5�1䌜;2�"�|�U��d��T�P����mBL+��TQ�m��
z��}�$m��D����f(�$�-Oq���F����y�$�����Qw%�c�[����CV-��®z�7�U3:1>�Ѣ�5S����S3��SS��a��L2X��NAlNO�=3����˳���Lc�Lmr<I*Q��.�S6�I�yj���n������"�EEl[� �Z�8dz�I�'=�ᰪف�d4��,c"��1M܇�w�-%�I*+�9"���In'�,�F�_U�dP/�(q�W+i�c�@��11�%�)�o�Sy�~`���	wN� 4���������F�&���'�dӦc���/b�����7|����+�7�,����o�?��'�|�!�� R����A���Oq�K�,[�p���m � �@j�������&���EI����������=3=��ȗ��V��X0�߻�����և�M�tjb2k�����}_��? �������+W�{4��>A]�S[��1��SO=�?���;�-[a����|�;xp|����_��ߜv�i�����@d<)0��y��ߏA.f\)��H\7��i��ds}}�3'Mg��>�h����PtX��t�pըE�Y�tyWw/F��j�߆����wz������	F��8��:��!�_��ծ]{�u���[i��(�b�g�\�<ޤ_
`��A�Zx�gA��j�2=�Q�m9z)�ر�H�S_n1��T5�H?�%'Q�����L��_�)��[!>!9�xC4ocH&�nyÕP
���.%�͙5Ń������w������"����H4oa��F��UE�KN��&w�!���+�#uY}2·�k�j�1�x��a�b�ޑ�	,8�.G��O�2�Mi?6�&>��� � ��ڴ���'H,�B��7\�L	�����HӨ� ��M��8��m�@��>���6#.� �[�]#s%�/J搞�B5�X���j����0��$�^$��Lh�7��F�[��!h�)�� �!^x�������?  pc���pF�̾���������Fފ7��o�R�+q��W��թ��
2���o~���g����&����~�G�	��g�9>>
nH'�	ya�>�� 5@���E�7Ρ�S�\���D�� {�1</��Ǧ�����������?�$�t%��I�0�T��71�������!��U�O|����k/��ҧ�~�����(�5���(�)Yq���/��R�x��1b���/�òe˞y晗^z�5��p�hO��Ѱe���%CC��Ǒ��yBK���a4ްo�S)lt���T�F�R:�9B-�+�#�Vg����6u�*�X�ԑq�z���g�5���Oװ��i�t��L?�P&Љ;wz�y��f��{{�(��r�W��t�:o�2��ņc�V;��7���2�̤M�0�1|Y��ݶ� D�L����I����-\80}`Wb���غu��@����:��ਝ�[ҵ�����}�\�8겦*�yT���g��q�ϟs�Ф�ȸ� n���4��`��͇���-AJm�V�YG!�1ʡ�a3�4��Jo�;T�+|��C9�y��ȼ�2"qݥ��,�yk��B�D��Б�0�r��#�8��s��ׯ߿w/t�əE����`�b)����ꀝ{�!놆������@2&��V��&���~�x�b�(�=�X|d_�b���SO����w�}���������׮Y���g?@������ �D?I�yi�A���S����� �30�%��,'�x�������)�>�ʐ��%rX�"�2h�R�]x���?��?��?У����o~����U�֬\�zdd�@�@V�Pc�Bb�������+�q����ַ������Fy~bN!�n��VT9Wp��я\�t��8rU]���>򑏠?�u0���:#yх�!e�a</�W�w�駟�s��n����`��|EԮ]� �0����L�QB7��*nz��'C�ɡ���܅��s�4�Ħ��rmsS���Y��%<�Q�i��YP<,���EͰ�&���4��d��yۮ?/�m5S����O�e��,��׆	*lT25��R8o6#�q<��e9©��|���:^�H]ԁ�Ya�1c�n���t�
h�Ƿo۶mp�
IY7�i�g��fzS&���X04Ȱ1�岞ݨGe��,������g�\u� L��q*A��r��=��Z�>�Kۚ?D?�^��<.i���&��:>��G�8E���j����@�]g�Rh��u�?�xZ'�x���������h���Ⅾ�7��`��ŕ�<� 7%����Nz�ɹ����O�8fyͪչ�bB��e�3K��5k�0��.���p���X�x(��Pxj+T7<�R�vpk<8��s}���ݥ�aw���Yh����S�����x�q�F����������1&� �ՙ��?��$M�"�f������d�ɥnv��'�B�n\��q�w��_���<�뮻�24.WHt�׿�5���{�F��>��3�p�ؙ �(?�|���z�Q[�U*��<Tɹ�}%��LdgA�0]��	���jZ��^։e��?�����f����e[�m�]�z�Io���>#�"�onZkT���\��v�<|�����-8�X�YkH�;���[�L<�hI����\4><j�M�gi=*K-�S��m6�jYZ�]�`���Ϊ隙�3 n�=3�EE%6Ugk��(]5��6�t���g��,q�Z�%�L�ԧ�k�N�5�u1�Q8���8	��-���"�m>�m����ي����%�+�<3���\�+M�'�sq�����\�M}�V�f>�e�ĝ����t�}���Y$�1�5�p9�jIe���Ur��q��Q�Z�%�ʀf ��?��?��7�q�-�b�Ϗ��oW�</h�X�fm!���G�c���]{���K�/<9E�
w�P��ؽ9�M�D=�z\ ѝw�9<<�<��R�>��:@�0%  R2Pcdb����%�l޼�� �y �v�_����}glv�],�T�UG���?9��?��[L��.�Yfj�*�9t���7;1>�B#S�s=�@��}�i��1��_k��X���>�n�-�q\v�9�S�p�qǏ_q���.Ϣ�����b/�Х������ecc#O�^% ��PHa�hN�d�tt�ndmɥ��@���j}rW<yD��P�k�US�c����Ħڮ4ƙVf�v�iZ��\MgD�����xoq�5�D�pU�[��oE Nl�+�P�`��ٯ�k�mYy�	~'��r�*���P�� 2$@$�$+Z�,�i��˫��3K�n{u�rϸ�Ӗ��da0H( ,� P"g(BUT�z��s�����o�������w���}��{����ogیB��@�Eo�z��1��e8�Ԣ��0ieC&���ׄV+�hh�,>����K�'yLRF_���@܃3�,�U>�(� 7��~!I���E/΅�-<T�ù���DQ�J($]`���a�h���Y@�+=���0Yyr�ؗ(��I��{B�V$�)��0	�Ex&��ݯs��31�#�|�{�We�!,��ꫯ�C�0��������P��	?c����[����v3!��߱o+�߬�O���񠥘�� -�D|����H����FEv�"U���xĹ����Ƽ��[p5!���\�'	b�����9��!F�'�An�a�z�P��]��-LZ�-�K��0ة�2����Mɋ}�:>��S�.A�x���T`�x2KK9;P;�Ek�-~�C��\��bVW3���uQ�P��m�C�``�T�8�L��ٕќv�9�w��Z���Ӈ����ע�9d��Ħ�<^Ą]F����]�3�+<����>t��_�4�t�V�7�m�V�V3�ٽO���n�י�� �ev뒩U�3[6�ܷo��d�j�-]159:���rm���+g�hr=Kj�J�)�]jo���2�VZ�oN���k},<HO���������
�,�j�~�ŉ�~���(+��g9�M~T���`e�\γQ�dmÊ!���2�fS|V\���aJg%f���D=���W��Nj����9ʺys�561>?/����U��6�)���{�G�VWG��G�:�Ng��~T���� Z9,ո����N%g����Gq����)�o����0sq�����a��[�s��FY�.��i�ר��S�}��I�V�Z�9�ngm��z ��( ZO�۫�!DN�/]"�#�!.#���SB*��ʐ*��ܜ��n�K�ܚo�y��j��Y�O�B�Uf�SɈ������@b$74ण���r��)�#Dqe��Wg���eX��e�
O�������*E�f(_�zc�%{Q9��zd�� �X2z�����3k�ox��ׇ\��8ߦ5���*��(�ٳ�>��r�ǱdRsT�|R�C-4�+-�D��*N�|M�z�v��g���䤐�B��ЖHEvV;��̔��:O-f	 ���;��CR��w����p#��Ԙ���r�V�!�v�����~G�ƍ,�D�zq�����>�����4���t�Ё1�4#ڱ���׫��1]+�y�	yt��V�^�"h��ѥY��1��r:\P�4�P�(AXZ��vd�s���39�{�V�K�Z�U+K���GR�5���=__PG�e&�i�#�7]ĕ�gi@�����)>�1"^f}+�;�-�$�M^���V�/��\��#L\�M���V�W��K�,�%�*@�8�!?g��*�nx��D��h��֛�K��u���@A�}&�Ny�/� !Ś�A���ѢmJH�$$��9*�@?��}bv;Yo͵��n��OKlr[Yk�\tn��#�>��hIJn�~)��6�Qr$�}�z8H{�}�u(��z�ʘ��o���>�:^�:�}�����-� T1B�N���+$�c�QL�W_x���OM���N �����[c�;.:V�J��R�
r�f�j�ϣ������%�`��\2��&�`<���-
W�4#�����!��R括���iF�^��n��l&��x0���.Z�) '*���(�u�
��B�6T�5�T��3:�,�T��TXw�E#��ϲN�����4��i��$V#KJI�=�4\�k�I˂�*<Z4�:�re�����1`�V��(�#obMj�ĉ+K/����A��C�E�-f�Z��n��+V�4�64� ���%�
��ܤ��ҥK)b߆�v����xJi���*Wf�5*" ���-;GC�L�N�i3@;���#|a� �%M.���#d��9N^��� ��P�2u{�ZoT}���2�\j�0t�t%�&O/H2��n�|�s��'F�-r�r>��E}�Q!��Ù�Z�zR�g����^�0t �������쬄un�.��W�^�O֭[�?w��������sBZ�8k�Et״wD삹�v�G#�aGv�D���on��87�R7/�P\ȗTB��ZQ9^T��;��h�j���	�ں�U�mɒ�~���,�r��X�>�.��$�__��\at�>=%��k/ݕ��+W���%*k����8.S��=6a����5����C���E�M�)�̓x��4���܋��SG��FB����2P�;&eL���]ĩ!�^.ܟ�:k5�=e<�R:Q��5��G��.Quk�4taX>.�eN�AJ�s1l�ٹs�du(~����>tSS�s ���$;B����I���j��#z��]�8�/:'{�G�.D�[���R*�H!N�
kBq4hv�8V�i���Z�l�广� B=@�8�H�f�M	yfi�}y���:
l��+H���X7�jG C����^餱�R�G���X�܊o�`8�T�Ͻ��f�B�#>Eq�ME�a9��8㳅�F�"���i%�~|W���jZ�	���Ǿ`V&L�6J)F"�+8��m۶=����<��Y����te�B%�|po��h��M-_�Իo��͛7��i��MN���IER��*@�R�=ɺ�����wχ7����
����ku�\�jd$����L�j)���^����:h�Z��5kVc|/��$��Q��Tn��S�F���s�J�%�ոݜ�޹c붝XӃ�h�+)�=&<:R����O���MV���6"3=%z˖�΄Y��F�z76�b��m����,<�d�Gy)3T����;�$���l%`'���v9Rټm�7޸aÆ˯�rZ%��.qE[��-[��կ��\|�����Kj�y�d�>2NK��j4�]��_����ۻw/}�W�x��?x�u�]��c�)3���g?ꗬ�V�����+�^|�^Z��i�|:~Qv�*���{ ���?���Kg>��O�MV�Zu衇V�J42�i�&|N%��ꍌ@"V�n�t�:�C����e�dD�4/ДD���r�yW{�EEi°��Ei����� �\����$N�&0>:�}׎={�P�.[��vv�����B��|)<h٧�`�bG_���6�d�Hq�V-1fX3�nҵ �7�g��c�`b�Y~LՈ}o3�!�-��r��r��y A����z���(ۧ��gf��a,�Q����[(%�Wb֯_���#�T��#�Q9���-XvH0�\l��#�8����>�9����D�՞��c���ii��j9�l�=]��LN������mK�:J�0��~�ɾk~�u�VP�����v�D��}ec>�X�%BY�b�,�y��ܷ/M�z����z��E&��&������%���!�k\8�3��v�d�n�/*χ^�Ƈ؃�m�A%$,%Jl�ow�.{5������AI��MrRqE+�$e��G>���i��XO]��O��'?����-0��۷c����_�?�x��@��(e�bc��/�;@d����O?���_��i5�=w�q�{��^\���K/��M��`��sH�RA4yA�;��JN����sN����n�\��w��gmٲ���{�[�^t�EX�_|�?���$��+�8��#S�s���<&��h:��lYD�����[�AI�U�3�xs?�����?����aT���O<�D�o.���p4u2F�X�dFpcs���/p�N;�4
�txF�/� �%.�W�����^ݱ'�U�Y6���m��Jз,	�,F����d�M��3	½�ųrr�(� 7���-�#Y�4`H`)���z�ꕫ@�=	�↤�r���Tv��ח,��J4˱��;��ǀ%��ر��<$1�mn^Z�(��"�P����~H��4-�6��4w(S��Yl��d�n�ɢj�onۃ��_>�i���@�dE&�
��W7o����A����o̕s^��@M<ߚʹDF(�ӆ��1?�O��+��=)A�0A�����m�Ȗ�uk,�š�������χ�<���o���\�$�+ϒ��H�������3��h��#��Զ�u�'E�Ǔj���/mڸ��k��Z�+�.��K?p����'F�67���.�� �`���˖-��_�����{��7���~��/%���W��i��`�����{��b ?��O�}bb�㎣����y��[jQ�QKu��6-F�������i����������w���?���΂�>����ַp����窫� �����_�K.�$P�Fڒ��jA�L�\���5�Y�I���e�u:��P��
������TE+��G9>2ʊ}PS�U�1TXF�Q�t��d{�9������O>Y,B]�R{z�fҀT���UE�y�K%~� s�aZ��h(J��ծ�� !,%�2�k���*�P���0mn���f�z>��w���2J��.��L���,�g|c�������"ϝκu� ��8��P+�+<����;����~��t�r�q��.B�6�q+�a��\p�g�y& �+V	�S���Yg?��c�<�ԃ>X�I��\[�x/3�:�+�Vt�d�����)�j���P�"�1h�����;��0�= ����q�~x&u�v�'��Ǐb_p�K�Y�����T��X5V���<q��5m��ͳ��ra��!�c�����,�^�m����e�u��b��b��� ���s�GT�ȇPg9#�7�l]�z5���[��Ē)hv3{��O�6F�ncK�h�M���k@��`d�(�c��o޼��ժU#����^���N:�.�W6o*_�z-����@.�Ko�g�Op�~�@�.�3,B�U/�'Nn.����"0t����7l�`)$8NxÈc|�o�>h�L��i|�W�<�L0w�s��7�9>1*��NY��f����4�C��7y�7H]Ʊ�>һC�O�\�f���SN�����y25�Z<K$��V�g1F���$�m/��b<˫�Z�_b���9�#�)Q�|��D�ȑ���kZ�i/����Fu. ȼ��]���_C�L)e��hyP��L���1�|����$������<��}���Cmӱ�EeIQ�I_�ѧ>��3�8cbl,��d	R9���W�\�?o���w6�%es��v�f����p�6�~=��{��qŸ`
~�;�0��O=*wHJ]MQ��������y>�)Ѝ����[��-Y�t`����	RK�d|��e�I��hL6K+�Jխ^���l+�jW��q�4ye=�.�(��e)R�5�n��NyvN��*�#"x�\Ku�DV򸈒y�����Y�T�^����R�S�A \�Bk`�~m�V�VYs��[o��������;�W����x���c8�/�����151	\y�!�K�δ���7^�w�߽�{p�	'�@m}���y�Ο���W�������h�vr%^>��OJtf��u۶o|�@"_r9��
��͉�1�T���T�t�c��e:2�=�;�̥�^
�I���~��'�z��kV�N|w衇�7��]s�5�L�����gIB��`НnK�)�(.ؓ��b��`�����>뤈� �?�0�-�=M`v<� t[�1� �_�q�Ee�2 �k�ƾ�ʋ/����S{1??+��$���Ͻ��G~ 
�ٹ|�rl�vފ�>�䓀�+V�����7���Dp)�x�ݻw�� v��u16��f[���\����77��4�vXx|�Q�}�v�-C8�xn��wsV���.2�(�u�|�� ����~��Q�������^q�g*"~}�kP��N��/�
�Cuö>��F�]	�IEt��?�x~v���.��%��pe��K/nz��͘Ԗ�^h�p�Q�s�@ڮ��xQip�3k���X�Y�_~�(��R?ddD]bs�,�}���b�mI������L�q��[��9/Z{Z�BvZ�S�j�Y.�v�o~{nF�v��~l� ��7��A^��p���x����[AL�QR���py�`v�4y�&�CX��5lc�����?��?��;�9�J���g>�������{,I�8���s�� </��"`=�)���?�8)
�������>��5~��N��Y�^LW���0�>@�h��"|����Qy���i�f�Ę�:�SO=l衇�?��p�X-(�ϒJ�=;G�j�BuZ<�̚~9��q�&'�@���K�|�>��_��{��b1ZN�[����&�:D_x��cRP�/��r��ġ`P�YQ�5�d�M7���(�_��_1 �賟�,��������k�� ���L��O|�rt����o�*�#������������$�7l�}�y��h&PxG"5 &IZ��{h�ȃ��"��0�r7��,����{�MiS���q^��'7<�C<��dZ�K�,�G����P�>��/H���_��UW]�3��cO`m!G��gAK�Yg�	��z�ǵf�4���@���w(�+.?��{����_������2~]����2p1Fc�s��B�K�I���NVz�I'���� ���ݤ�s[6��س{��,�i�l��nr�c+�W^�^4㼗�ʣl,_Um��I��ԋ\�E��H�4Υ�s����xH�uq�uٳ����8�w�;W�{Eu,���H���z3�@����Y[ö*ĳ![7��-�ާ�~�4��z>P(1���e�YA����:�v3v�*0�)�y�N;�r� Y�y�]͠�{v�>�0�5����ؓ��n�(���^�vu�9319v����+F��dMu6譖MNy����?��@�WkT9��s�w������O;1�8��b���ݼi_(���?X��W_�oN7[3�Z	+�hL�P�I V�M�U�p�\���g�c���s��̊�+�
_y�+>t�/��}�0�j]��{�4���I�����G{���=�{��ݱ����s>{��h]L4� q�6�LJ�`�+պ��^JzgVT��.�����;�~�ӟ���j{�de���X郗^����;�cǶ��;�d>��ï��JM��p�;Yg��������9���,�/����9�+z��-a���彧����~���/���O9���6����(-�����=���8�#��M�@f��i->��Cw����-دLjVc�#�oz�I�^9��s����裏fL1�O"�g��a�ȩ�i��uq@kL�-��
������`�id[�S�	��!K%�SQ�[_f~����VAa+�"���@�WWD�4�X���4�;d�Cܜ�������f��۶������q�v��瞛�� @Y�z���t�%�^0�B�as:8 ��֮śg��112�|�=�t�(��&Gv�����m�m{mǾ��yփ?2�u����A�ӾQ�v�XX��]|�|��u��%>�b�>b�>�-G`��;F���4(kj��h��؉��i���,��c �T]�XE�ֳ$�F�#>�f/)|&R ��Í	�vxMȠ��@�E_�
�A��H)�����0���B�9ׇ_��烑��aa_�E���N:	mH2f�e�
��iy����-�LzD%R���I"��G��qk�:+o�j�O<q�a�]x�|�T�R# s�����'�d�� �}˷�|�\s
p�����~`o�M2����L�Y >`��9�c�p��yfW\�W>������ukD�>z�eֽ��_+�%	N&�)t�O~� _����^����/���q$� �$�Ve�W��p�{�z��WK�wf��L:�я~E�ݹ�h��;`�N8���➸	P9�drr��{^p��eI�q�?C�Bm	���y��j�������_�+t&h	X
�<����6r�Q����b��3���^Y�إߦ�X3�s��{���	2��Q�@���F��^xZ�a��X�|9&�^�UP�5Ù��8�w;Uj׭[���d��%�tť)v�ں{7���rlq+���g����i.kY=qH{�r��	~��Fꢶ�f�RN����d�Ӟ�Ī4��ڒ�	�֢��8%0�.�w��fvv�9��w<��8IU�E��-S�Rc�A,=��fHb?노VFG�[��h%�Zډ�f��b4ت�e������(x����0�J��H�t��~˹�x}1hl�|�J��o �zR7NQN�8��8��n�Km��b�7xT9�ߚ�m�f�#{�Lo|��j<ܧ��sV��bO[���c6 ��:����pg�*|�� S�n���^���h7��E@(�conي�C��w�/���˰mێ\#Aiie���vR���9h�P�1�#7}��|�cs]�#���?��O�"���L,Lِ ?)�T��ٳ��h�W�4+�l�&����g�R���L�.D,�V��Mi'�G�J|\����u��3�qӦM���*���o��=���p�y}1L�;��X[����{�����^B��={hǨ�-L3����q�!=����1��3�P�
os�'��k>z�29i�"���e�#��q���!I�^�[I0�/8a�wς�'��&*�gcn��L"��7�I�Xfy��X-������@�̞�f���GNg �����	��M��A�?����q�y��ƹc�Yx�JK}��B)8�z��ږL�1X�B͂��$$���Cȥ��
呾rr�CyZN��V!�	=��I.�R=����fR�K|�p׋A�T1h��8�����c�.|�[`1�/y���`��B4:Kᅸ���s�<r�ȉ����Kba@Bx����뱪�h�v���Z���_��נ�}�S����s���\�
�O��O
��F;#C�j����n�k������8X���ފO�� ��?�0P�w����}w�{f|p�<���Ν�n�ᮻ�­p��vA9��Ӆ��D����kEb� R@Q��կ r�M	DY�|	p�UW]��Q�f&�$~	 �£q~�~�Y]������6l��뵺�'�O>��������+V,Q�J���Y*����L�ᴘ��a[qu��~�_x�Ygb=���+�4<���w�!�������|�o�f�}L
������A� ����x:�<>Ĳ䒝4��	3��M}�+F���,i���w�؁�c����_|K͐j�{{���l����D>�f���y�Аlb�'�}^n1؉р�k�+F��g�� �E"q��m��?�056}? �MW<�1?�#��c��u����`B��	�;��GE�d�l�P���:�Փ��(�T�J���,�Fl���f ��i$m�S�S�z�\������[�ֳ"JiM�\~�j��iηW�X��tI�V�7Z��^��N�^M%�R�\d�"�y��Ut�#�P����qg[kqdQ�-�[�Z�}��p��ǿ �/Z`�r��|��+�i��sln0�_8����[�JZS���C���1S;~�:m���iw�p����ĸ\��������ל���&1D�P̳��K����/��-2�V�f��&�'�����S$�~���0�L��MA6�z5x�Z�ڵ��p�Y��Gj���f���_����SN9��Oϵ����*4����;��0��/z�|�%%R\H���es]��A����ˠ]j%e
Q�t��%�V��a^��'�����s�������}211��}`��/ru�ϝ��������s���<�ԗeˤ����<�Lp��������1l����8�Xd̋����o�˿���K&&�����n��ƍ����_�~$t�}�#x����ClC�n�펏}�c�Y����~��nĀ1���>�������[��go��{��7���k�:j����|���1�/��w��}�������o}<��CA�~��gM�VRZ���8�"y�{�
o����M8E��M��+_P]�yUҌ��m-Tܽ%���|("�1�Sv	]��c��pj��1�x=x7���ć����r_��%Y�c �?�P�6VQ=���Pܪ:2��V>3�/�{���ѿ��~�V�ל��D?���ȥWm��  ��IDATvV�u�ן5d�g�v�vp���7���W|stF�gUkG���G��2D䪓���og	�[�#��ɾ�#��!���wɲn�P��=��;�J�x�f��pgfA?eց�RP��� %u����T�,�v6`m2W�A�֣D�� �SO=�D�'���o:���<i~�J��Xy�C�E�<��HsOS*3�|�K_b�5��%M�cZH'L���g>c	u�V�к��!/z����uSvP�LE{��8�(b|O��ڹ���]���]{�~$j�R�#��D�� �Jl������zm��ꫯ�)�� �97X9Fȡ�L�c�`�8�G}4�8�<餓��Y���# 9����c��o�&Bd���[�,�����z��3����"�V��cx��:�S֬Y��c}0�O�ٯ��@�dl{��ӍH
��q��.}g�b�;+�q0n�s�Ν*��;���ڿBac�������8��?�я�����q ��2�y���o�}��Ƭ��n��+G�o�D��zzZr#�]h����Fp��o���cI(@�&��s�$�9�j��W��+��N/���r�*��=���#�/�����_�n���>�SZɁi��{[�n�
!�8ɢ����z⢊nm\��|EG܍�d.�"飱t|��x�^��A/mK+���x�ػ󉈆�m�g�?�-~'X�_@�ǰ|PU��vTtI�L����tFX�K=��Jki�������͞��N�[�M�n1;?�f����&]u�j��v�	���2����������N92��g}T��K�L�j5м��Y$�X���
\�񀽓B$����8.���iݣ����^�ן2��)����rYS�a'-�yW8X�Z]��N�cE�,���c��|{>CHJC$�×/_J�d=�/�0���/��Ӌs�c��>:r�1���Y>:ƃ3?#�u��N>��c��6A'��D��ɲ����W@SSK/��Rz�|�e�������C�I�5t0#�K�2~v������n^ nh�{߅���Z������+S:�Va-F��Ptǜ��4�ng-c�.��oӣ�3dm�!<b��ϕR�d��:uC�5��j���l��]�&]��C��z�ctK J����>�����Y��_�!H}���8�@��ѐ5���ԒI�i6i�����U+	����M}���4ho.�,�ɻ�����AL�e��ҥK!�w�4!����_����7��%�c��E��&��Y�Wb�+��+ ��l�_3�֜������m��G�w_�9�,K�����+dك�[^�O<#ܳ\�ȗcu�=Gd�8�O��U*�ghG�PW�B��1gD�i�=e�̊�C��8����`� �r�BZ1h��h�䀙�H��ƃd��GF@k)%�E}�V�.�q茏��q[x	{1s �CR߆EԈ22>�+���ꪊ����+Y�|����V)�n(�����ڤ��P<�5�=�)�q��cv�g�܊M/٤&�i�t�Qm��R��ש-�B)-WTAX��kE�M�bz(&#���+2g���P@��8�R!��,�|�a�;{	�DA7�����J���>+5z#D�`;eQP*�_S��=�������_�Bwe�9�2 K�iӦn��q�y灃�eg�� ���?�����G���$;�?g��k��o.��|&L��yv̚�n�����AP�$�/ʵ����ץ�K ����n�1�p2?�{�9;>��u[�5+Wd�4���e���+�Jurź2��l~��<9v0³!H����n�ݢ�9!ⴒI�++��{E֍�^%*zP��g]�V+I%��TA9�@�s���{S[���k�K췃�r+�Q�G�CI�YVbo��W�0l����>+ĭ���\|�)��s��	_��n�Z���y��^Y6�O�*Y�z*H�n�/x��R�#{"ih��(�ki�<"�!w���FV.�>=�5�z}D���:\��i����}�#/�a)cu��r�n����D��^^��ĥ�라���sߐ�����Jt�blX���)6H�my���Z]�uی0� �'�2����vS.@�X��"M�g�Է,)|/�)ӹ��,�����f�8���B�:b�$��(@cq!�qR�6@�:�q��ݞP� �����R�U���J�Mo$�s��Q�-δ�*��U�����|W�z*k����r(�HIWy��3y�¿Ei�(<�g�/H28prUDc��g�;�&9B8�i�����������?)W>��s��w����V�0�F�Q��;BiV����:���駟β�t,_w�u����3Q+�d�Ҕ\E*~.����u仒�Y�[:)5!�֯_�I��<�̡���K�����u�|Q��굵�51r�y�z�S'T�����T�(�,��@��&B]��9�`��{��-^���a��ֻ����|ƣ�E�3_�?
z�vku}��cC��_�̠M�۾8E�o�!v�4����� �(x��w�3�y3e	�������wG����J����B��;�W:�s�Lt��,��ˉ#p}|W�U�y���`��<�3�4����y���p&2�ܷn"?be�^�l{O�q���2�׀^��-�[&�؇d��"w.���R�W���N�Et� ��DD.����l%)�y=���e�;đ����g8nC�f~qAw'�,J8�=�~��xx����\���A=d~+�������M�|�����wXd�w�w�E�3��K"ѭ)mq��Q�� ����߃A�'�����7��I\�'��;J��������A���Qo��޳��͖/_�Kkz!��:{�싋�Kk�"o�َ7�Vd�f#�x+r���u�T���;��n�]��jw��̼SD�D0Dn��l��׷��a���[%�f=��P���Ι�\��C�
9����[�k�^���3Mq�B`ϊ"�0fj�e�ەF�^�$ɩ4�Ei.��*�[��8lI���X�YE��Y�ZZ����F.��s�����w���mK7�cz�f84�Z-N�e�e>��b�q���"��,����q��W+4�>��*&0�!��V�r�h�p������3I���&Vc�S�VL�R�M��e�M6GB�P��U�)���a ���r�R�I��V�0��y\BT��������B�p���^h�ڴ���������d月��6l�����m�c�R��q0>B�4r��`|H4h���%a�@?�Т ������4��,�,�.�}x��&���FZ����b��%���6���׹d�H�W��| ���c���2���D&����{�m����:�^��s&����6!L��(�VՍ,\bb���ս��RQ��������~�{��O�g7�����X.�>Ჹ�V�/z�Y���]�	OI���9IIq�'���䏙Ӭ_?o[[�������o1hD�}HlOaQ�C���Ar�FQa^R.(�F��<�"_ν�44[��q�5��(.���P�������N�"0���%"Y��l�&�^T�|�i׷}q}���JQ����4�4׶,�o���2�Ƅ�Q�c�"�zi{�!�Ne�}�y���,�wK�r�+��d�k{J�V�,+��8��ѝ�!fg�,RM�x_����0��ca�EP	��So5`q6\l`"<M���Ł���x�[��r�?�?��/f2	j��-�{\���e����Kʑ�$}Y�{c-���{��m�=���H�j�봶�n������|�[K���ήn{E��5��nQ�防�����\.{&�|�u��z�9:VsQ/J��<�wr����*�ǽX<B���n�t��δFݞnkbb2*�V����E��Ym���&�����E�4�� W��x1���$DU�=.#G%���Z�F�
8���*�KÜ1hF��.�����J��iŉs��V�#$����b�i:�W7�#6�<ri%e9�"zI�:���3.��ڕJF��<�X�������D;�&0��?B���_�&�<癯a���)�Q^�
ןf�6F"7��He�s��X��,�LY����GG�^fr�X��vH��e���m�=_ٕ�U�K�?B
���/�;���LH*kK��.�E�Q�]y�1u�X�3��T�M��C��?����e�,J萹S�pt��w���@��h���Ow�7*�ⴥ�y'�U�}� ,�N9dV,�(����m�J��Z_*1װ�E޳ϫ	1Y'�-|��*'e���4i!{7��;���<{��U{�Qg�]��p��!��ë#�1���2��x{d�&(F�����R�"Wky��VVoHHI}f�-��U���Pl��XvxY�:�ǯ�����Ǉ���ϡ�PKYh�=��y���{L�����yE`�3ǋSNϕ0\�H��iε�Xe��G�ƾ��~v�G����R�����cN3���׆6%dE�hx0,�Z$羐[<}W�v|���}}ח{�J��b��VO6G���
̔k�	um?H®o�w�d�	��Vɕ��BkO��zã-ϋIYC覧F�@&N�i�����MH�h�����N��MR�D�O�k�1��b�E?�2/���V;
�%�����bfZp ���N�5���$L�����E��s�jxq`��:�1�7�~��r^|�Ы�Yc.����)�k��n��	ЖGf�Y�m.Y>!eT!V�t�4L���)ґ��ʞ=�ذ�zћ��v�;-|�1���W�y��$B8o�Q�5���Zy����Zn-�S$��S�.�h���,�3#�z�'��?����Q,���z�s[�pA��V�f�i��5P�훗�m3Ժ0\W� ��0����IDZ\H$Aq���W�ޑ��}�Y��l� C1B7�y��P�϶zk!YT5>�j�@���[U�S�F9��8��������3��n.c��7��ϳ� ����?мj<ϐ�J��R�X=".|[t���C�#��KV����l���oŶ=)XFw�	�жڎȶ
}��f�'{59���2(�٬=��,;<Z�>�r��Qlnnh��(����߬���&��͎g4S��/μ�qiRH�N!v����|���oTC�/�_F���W� �;ltE��ݤI�l�yY�Wx�Dus���8�����M|ѕ"���B���/�!�u�ε������e�*zu��;v��DɊ+�bf�<k\��S3vtt4���V[�~�RE���y����h���&oڈ�����?�=��� {Q�O�9��������b�GJ�.�Q`�s�<{2껕�;N���g8�f_#DK!�}� 9��2���9
�Č��YÇ�EQ,"�8�������D�,�OT��!���zUv}�Z�!���n�w+w���-�e�,^"�� bMҪ�0J��<�`ֺ;F��љ��Q�J��zJ���qR��	i� j����/�ħ�:�ЋÑ�7���NC��>�&���|?Oy�ǭ�U�����ׁ�rZ=ާ���gl4�5�2��	���l�C��)[R� ֋�knZ�\����:-N=-���d�[1hK)a� ����ڌ6FXuw�޻�[�yzGi�B�4$H��A|���5�1�v�ݳ}n_���\%�ӽ�[Ŭ.zYg�X�t��d��$��&�kT��(.���NO�z�7W�:dfVR��ib��&��mI�´^H�+ ����ZO�N�L��lHy������9Px��EyZ�� �Z,�B��.7.f;�*���ڎ=��<"�YF!(=:��z�����D)@t���.wWu����*�O��`ez.�'�����ؙ�V�5eM�S��5^��;�.�!*���\�\��ڵ�DXc)FQ���N���r �S_��8�Z`���|���^EM1-V󠢀7���^{�6B�,�,)�8�i۠L�����t;����ݛo�	a/ͳ���%c�9�~��k
o��]�<�i�B>"}L"q��ݦj��x;) ��w�L쉽��B��'���&�/��NAOJ�`��7.~Ҹ�mk3�2[vE�I����@#I�MW��eU<������OW�i�e%t�z,c|�LR�����3���Kq�����()�.�Tj�nY�5�{ʏ�����ä�Ny�����E23�=�\��d�E���\���4��)ď��'��
��p�r�q�f��:����0|��iB�^�z�r��:6"u?�=�e�7�lٲu�6���FO�2�%(��BE�׺׮_�>��333�z(�p��Om߾�КH�wԼ�Z�8���2�I�� k~{|��Y��C�ދ.�:K���,$����^}��];{Guԫ{��&H���M�W�\)c�E������4R�~�us)���+	��Bbkj��9`gxDWyH��+d�6�"?p�	�x�\���/������'�b�ܛ/�B9�
H�\�4��i)��hZ6��y�����)z��s�s�s��m0� L|Ec ]q����[�C��=�lib@3nx�U�u��M��KuM�kz�؜!JJ8Z0��H-u�!�1 h.�:Z�,_'�B�q���{eְs��gʊ��0F��V�Q�}%`,�ᖐ�bF��|���X���A��h0X�P�O�	k��F7(	ث~�\��FG�o4$
�e�z��9���z�b>�@~�n읐��j�(DπR��S A4�_������"���V;UU�H)�^{�5I�VC�5.8`�j����۶m�|�$�6�ZT��9�ۢ�)?��3��,�]m�tR�m��Iq��9q%��\�r���S��̛3��|w.k�ϵ�X,Y��V��5�p|b|)����8����|��o�ܵs��b����<��C�m�*Sr	�G7K�ÞSYO�v"�����jL|�������b|+��2�n��IG��:V7�$�mq������>��v*4����va�U��/���Z�j�*<�O4��u&�YrL�8�`�l��n�ب�K_�o���Rw'�b<�4��?��=�c3�ʙ�kx7��	�mȪ�nb`Y�w��g�b�9O��M���L�JY�Rp&�"�''��&YW��/fWo�j�����Z��t�T�J�����zf`�e�9���Ͳ29m��Q@�eYD��}��I�"(ԕ�	�g}Dv�nr��dJ���|��N�ZZ (P���ɂ�u��J%:g{�o�Ű�8.�u�s��K	��Y���!qص��Y�(߭W�Jr�!I�K���1W�28K�!a���N�s�
[�*|�ʈ.u��%�etM^�!�0��.0v���$��S��if�h�"���.�C pd�۪�V� �PæM��M˖-0ݷoXN�R�o5	k�-�=�.]*U�gp�?�tji,cК��"�j��x�������D3̯�C��E (��L�w��㤦2B,c>��4��J%*�ha�#_m�97�1;Y���=��T��Nś��q�?�~�B�Zc,�^C��^��݅,����N���V�!Xm�*
�b��V�ŀY���H�c`�Na��RCB�Y��4p���V���E�2����G�y�I�d���D>r""�8�y't�ݨ>��2	{8�>=���W��z��=���DAQR��/<���=���ed R��:}`�5C$N4��E�Pc$1�ݸ��J1�����x���x!�bN��N��V�6��J�"1�������ȇ�E���m���AQrC���y���\3;3��w�ցт��@��1���~���	ϱss���eg�/�j\)�3F{���^�}���q[r�G>|�)�7����Yr6`�3�<�SN��Y��7��̓mܸq�֭�7o^�������im�S/	�Ǆ��{��ּ����9�s����橧�z�GQA�E���EF���b`�^w�d�u>:�xŊ5��ɳh���T����FG�fg$�tϾY n�@}ϴ���fc�V��kd\m�vW�j*+�$��YW,�I�aع��*�uI Q�I���8/��:�^�p�~����+�C'�Xh��G䊝#�
�J��#�!�s-�7���0(�=�HV�\��f���Jjf"��T��IUʭH{ �uqbJ��#�,�;## �]����q-�=L�[�K��8��W�n����DZ'(&+DZ8t_����&,y7<ET��U%WÆ߻W���jU	��Y�I��;"M�m����c>��u�yF�^��#OƱq��f�
�᰽Ґ������"��%�q�j�uRe�1�g��?4�pY��Y7�-���ܓHS��C-�c"Y"m�N�K�Q��Lѳ�|��tJ2E�+$E�*���zkLi�a�\]p��b�`ʜ�ZE2Z���'�a&��2�^lأH	W>��j�+e��8.őиOL�@C��}����:or1��?$�\#�Y}��@�PKA*��Y*#fy
��X����Q��ݟ�~�y�Y�=餓>��O{�p���<or��G�qg�}��~����{���&땨S`���u�>��1����v�����SO=��C���|����p�����a�v�m�n~��H�4[��ڻ��\-�>��)���$1⸪�i'�4==�]l(F�^��t���^�X�N Kt���N[������-?��}��,@�ď��E�gm���ʐ��xAU������~������o&]��:aŗ�s���|�W��i�3�7�x#�0D=O&�������jV�^��+��摍6lXw�Z�8�qϑ����O>�$>9��YV�ꠒ�s����k?��Ӈv�����|l֡	h��+琛���h���z}��t»i䍂���u��P�)�4���>��h�E��f�ǒLd4fuA��nC������Ҳk�9O{7��z�,�B������E<M]S��`(H��tRߐGSOb��0#���� pg�=��#������~�L�!�'E������M[�D�-�&��CxǓ�6`C�Y&T� o�õ�-�-�P����G���|������`ʛ��7���:��?�=�y��|��G�"T�8Ԋ���^|�ŗ_~����_{�_~��W^�S�Ҩ&n��G��h�62jǼ�g���7���b̔�1�;.�y�3]�jZ{���^�j�ڔq=���ݻZ�nkY���X#���ZMHC3��$��Q%�_�j�`_I�We&Ny�T�n���'�c �Ӥ
$"ye.:"(<�T�2wh�C����.��u�>�����6/���Ē6�\㒥=�z����D�&����V��%�Vh�I�U	4k�葏R��~9S�U��<��7���|��wNM�\$��:G�{D�8�8��]w������;h�z`S�|@8b<�Yj������o_�v-g[�u�ku�K`��Iq���{������1����%J�w�0������X�E�_��:�\3�s�������`y��ۿ�v�A�|R(w�����/��o~���K/�{��oU/_�;�&�?���1��~���X�vy��=�أg˖-w�u�p�	'�6g}�O��k0>(�����q��x���?||T�}L$C&��N�%T#���z����X	��NH�C�5.�H�\�+ܕB]��P&Ra� $�aN����dI��jiVR�n�$_�j���^�͹�N��NE���F&yO5��EI~�د��D����"�R�&xh0윦&i�/����?����E�J^�6Ҥb�#��G!�ɭ���w_{衇(#!w�?��k���j��6m��H���^�>�NC�`�g�u�e�\�tRr	�Nv�؆���Ͼ��K<��.��Ï<����ʞ���:��J���2�/j��׻���ZҺ�n��k5�{���kr U@3���i�J�Z�b��8Lw�C>\�B8/�U#�ܡh
�fo�H�H�v_+�|� E��A.�g��s��
�k�:������B�b��T2�����3_W��$)S�}M���4�F)�m4,1c(o[u�r���7���ǩc)}�Y���$�_����o��_v�e`��/Veu��6¶}����{�=����Nr̶�o������w܁;����mb��9�� ���ۿc���>.�Gpe�zY�B��M7��W��t�kVW'_��z�\I�t��}�{��i�jƵ3BK��g?������ ]q�N�R�O��}��5����$���?�*�f����ձi��8����s��SN9�\�2�eY�R�,|X�}��������Ǿ��/B���˺.�MF��H��������XP�R�|����ݿ�w�Ї>��OiK�9�L��fI�jV*e-�y�M7|�� �11<:�2Q�����n£/���Ls��v[RcX�'����{���,;_,׶rǎ�;�|oP®]�~��;��Ɉ^w�H��C� >��C_|�E���2d����1�3Π��zff�`۶m�V*ƒb�V,_	ٿn�:���~��0ϭ��6�@�a|HɆ��s�Y1>:2�hg(�m��æ�����cӳ3�؈��yc41&͛Gj��;�l��K��h��F��E�"{����Z%����Kz\���+�K0��4�qR?-�c)B��;q^�U;��
��(�d9K"y�bڇ�����
�eI�Q�R�#�����.}�Rc��pW g��z��,!�'�$J5y����c�(}Z� Mhb*�-�ċ��֭�ss��������F�\X�x��H(4�u;��Ͻ�f������!��b�
��,�H}t~~��:.5�����SO�"�i�[�LX���T��{��G!��b�EetG�C5|�M�f�P$���C�N�u�d�N&q)i^���O�3�V�Z�#"��-| 5V�C�_�����QGE�&bAp��b;�^_�.����Sm�����ªdd�.� Kũ��u���16���v��G���?ICka�����y�����X�t��εS˦���W�������|��;���<�@ZB�Βx��=j�{t $b/ڲe����߁e���R:*0���A|��i�T�K|$Xv�w5���1�U�Ș���B��z�b���:yF��>T�*��g3_oV����}_?�+ԏ��U۠�$�V4�CX�|��4��s�=[�n=���G8�,���Ѐ�c�֬=p��=�q3�5�8�D�gAa���&X:(tZ���9��añ�n�Ï��Y<n��p�"�ɝ�a��!{��8xWj�Ҭo�n��3\8i{~F	@S�F��G��az*|Ҋf��9���ڷ)+��;YG�j=���n��?��k���;��9%M�dY�G���;m��.�F�nKS�漬X���n��@�Coo-��7���"�_���l��o���t�A"ػ"��A����ǳ@��^{-nf��:r��e�6�	�=R����Tr�g7�m��~�b^Ɛt����w�}7������_�~Ϟ}���J����qM�"1; q@T�
:)}�>��x�1�pnܸ��q,ٲ��9)�/����xX$t �~���d�mK��k�-�����͛W�^�������I���6���?�<��G?�Q��=���%U����.�ò�x�4�(#�E��Ump�oAFB�^}����B^�0I�� ���M/c�ps��;�)p��G�q��n����O|�e��0=+�)�~�f�����c=Ǿ�����MeL�	~�T��9<kƲ���~�w�)���d��L~]�,e��d�w�F����b�,�HR�d$6D�>��	�$�:�w>�������{�9��[i�r>�}h���Ҳ�����5���մ� $f�j
�g���<9�	N��e���[g�5<���w�I�u��/]7�����#�ՊuN�K]����p���Wc��Nǵ�B�J�U�)����°�@��N!�F��_�C�ϝ�"�K��1���3�#���3�� ��H���|�mƼ�3���E-�(�ۅ�7��ڱ�<{��Cw���m���Ō�M��I�\�T�������wء�~���$���lQZ�ˢ"�cc Z���s��?�C%	+�(ƙZnGN`�	�x��Z��٨� ���iu4�WUǖ���ن�`�ѷ^_V2�I�r˞��o~�x"xA�Ey��a�,���_��-��r�YgA0 ޲�2�pH;���>��������f�J�����o�5}�����S\������ɧ뀳���o�}�ӟ��8�`
4�PI"���Ï�b0����g�=11�x�����WP�`���^��y� R��n3;?;��ex�n.Y�l�����l�;���W|����ص}���K�D��B74���"z�-c�W\�!�LS���R�rh���g���_��`d��%oɊ��H�ʙ$)0�!�ʈ*�W���˧��S9ĩ�w�-:�� vn14	�[� �A��mݺu��|�K���\����h5��V��%��N�6����x�V���h6E��]�I��Z��_~��4�����׭�1ٺmg��=2>&�Z����%�z�c�ӡ����f	�<��b��&�@1[�B�Hجjgj<�� wL�f�~|�(�u�R_٫P����4H{9�0a�>Ý؟Ե���3R��Y}η��s���/LG��7�""�2�<�v�)~A�6qB?��> '�t*����Ж(��lLMM5`P��;��_�\��9n+Muq��
-��_�"�A9֊o�D�g�;��Y}���'�K*eʼA�D;50��)�K_��8_sY��q�e�w��~�~���/��e�Q�������cM�������fn&u�7b$�U���.���+����ӝn�G���5���c��8��M�Yyd�4�~��N8��ӱ\�!�ee}Y���Bc�7�t����$N�ωW|�8����C����կBr ��J��".0ˬĥD�o��o����韎<�H!��u������>�l5���
� �D����{0Z3D���|�k_�WT'��g\�@W�0�a[h���}��Km�Ȑl�c����Kl߾[o��O��OAҸ�3O=���/k!3V+s�ᇿ��~�|>§��9zE_��<P4-������Tz�[��ƘEv>��N������N����ݶc׫��1�w��Dm��+��0���T�
��#6�FG*0]���ϊZ���:Y�6�e�K[�m����DRr�+��c�@�.ыSZ�\�Y�
���J�<γH���gs�=�N!��YQ��y��om�^��i;Z=������mx�Ԓ�(���9	�HҲ�B<af�N��Ͽ�{QySH�Mڐ$l(���'��x �^�71:�h����+�T֞V�z��j�ܶ}rl��U�[s��J n������77V�U ]�ǐ���iq��O��|�#���];!-p J#]^:T�H��lA�pOr&[A.�́�Ǎ3�ZD$Ă�k�b:���,���t	A���(�2��+�5 2߾Ҍl���#w�x�-����WM��~]iU����D�`�zX*(����}8���>�9�kl��
9ɛ�)!kb��%��SN��?�=�H�1��~�$��`���j��[#c��V,�7��W.���N.�*|�;���Z�ob|�֨s���G�d��e����$��2G�˂o�������߁�F�O��V�Ů��S��k�-[���/u�Q�?ʝW���gd�&~h���D�L'-Ou��g�E�2�^C�;
����F򠾀'�OO<�D�|V�y��j�#7���>�0:Z���+1�Y�A�P=�9�,��/�֭�'�q-f't�]����O<�==EP���8��/|M����+&%h�:RjmZ�Ej�l��&6��gؘ��W`@on���]�}��<��*R�?���X�����t��Vv��i��)���С�|����e��V�ﲡ!E����z�yIP�����|ԧ>��n�r�Jh�@_��W�̤����m`�ĕ�/�ƍ��^t�E�KZ�����Q��%eC�=���;��M��� �m�d<�1(�����3� ����=�!�lTĿ�Y<� *����.�v�{ϐL��g�ț���M?��Ӏ3�{,���͙�0�α/-�����=�\|N{n���}�!N ��B��J�V�U-|�C��~��p=�G� ��KzԳ���a��z��h�<h�j�n���pA�Y���ͷ�g��kX7>��IEV�K�U�G8�'0�)���0_�ޤӞEv�/�of:�uE��6��10/	dX�bx�޼��b(O����g�}Ș��Z;PCzm�O/��J�X�	���{/	{��޻�˽��0k�)x8)�>��TO�5�@�i�"bx�G��C7�Y~�j��������Rղ���&���<�������K�,��2ߡn�-'��(J�J�^�e�fwllj�5����Z���{��*Ԁ"��q��W9΋4�;��0�e��#���Jd�릮� �%m�B���4�g�>]�������Еe)�fJ�y�)D�J+��+��Z�k��"����A��c���W�Rjw�7f����� ��K�� �#K��nw�� ��F���?�``:�އ���n�A÷o���xs��f�%)J	&f�/�?_|���o���~��Y�R�Q����_��������+�8�s�n.y�(��![㈴�E
���op�O��O��#_����[k�k��a ~
t��,S_��"70Z���������֌}�}&x��*������E���8���77�����C=���]vfa��|R���vQ CFBa�ݾ��/�ZHы5�L�UbF�Ej��`��r�'>��;�h��G	��v�4Ι�����L���JMd9W�� t62����{��1Y�k]�%N(-��D��=���K/�0�U�h/mw;DɆ�IBZ�Ғ�Mj-#P-q�S>��@�������i�"I�>���Ё��z�jȕ#�>J!�@ɩ%��~��_���/n���k��6(���ⴌ��e@<�r�O=���N?'�a����ǲ��Z���ΟIAA��H������{O� ��ڥ;�Ŕ�ai���
�ā�{�`�Q��<�&����vy�����9��tDB��F�Fm��%_�
���⭯|��ū���ț}m�T<���G��y�V�m���K�`/���zP�UW]ET�e%@���R�U�%u~��V�w-��,�<!]�?��v�mGy$tF�!�B�l�UI�x���SS�M��F����/�̓��`�Z*�]�O>�$DFb��6��t{e�w<����E*�l``'����� �}�"�-H|Q�c����j=���:زt�/���[� y#=�Y�Ԍu���_���Z��q�Z�2Ɯa�G^x!�$�	q�Zza�,��G�!ƾ��/�����@H�q�%K��M7�<x�1����7M
���<�r�G���\r	�5�5c�0PaYa�'�����ܽ�O��O!!�vzTD���h��"�rm�"1�G{v�8_�o��dзz9�-:_M02�+s�.�� ��,�ݹk7D�?�õ�>��Ԕ�"'q��B���k$��	��;V�Z>������/��[����w�4?�5�E�\�5�Kf�.�C� ���>�m��N�kH͐ٹ�������/mL<�س#���������ĊNR�>�z�u��j�,O�γ�Հ��ɊK��H-o��p�3a(튜�$���1��f�����o��ƮYA�ص�|�9KL&�V����7����Ϲ���f�T�,ɒ-��'lc0xbO���C�@:��JVH�W֗�z}�����[�
4�!	���b�1��۲1�<	I�5W�J5���{z��;g��^����*�޻��3��o�lζ��&�c�1�IF��X�*ex��2T3�]�D�KL�3 +�:)s�2�tvܤ(a���Β�Fj;�n'p'6F��5�F3��2n�p)��餤�t���}ӛ�|�EX�\g�<l�˭�Ep�_A��#o��/lߵgק���4���9^ƌ5��p�K��#WM	I��G��O��#�G(R��B�h۰Q2s�y�����M~��Ë����_����@�lnna�Zo.,�luE�W�M�4	�����߉w������8☿�D�����F��o�����/�+Za���X��\L�ժ��!���}�{�]w���_�	�����&���t��W*��|����VY��`|�N�̑�St ��O<��C=D2��9P�o��J�!FI��͎*l>6�E�#J#=2:DC���!�z٥��{��3S3YV����)��i7�� K�&�J����7U�
�3��M3��GZ��� �an����ѕCõJ��H��@��@��C�β:x�V�������zM��.�ZRM�-=��B����K���w��j�+W�P�K&f؋�!�13I��/�~2l`D�A$5U[�n�Zq� *=Gz�M0p�IM�^����&)�������7�.��RZ����ݻw�|ڱc��Bk�^���U�N�_�!Y��*�6[1�̶��?�-ņ������!���_��Ž���Q.���8�1�8:�WI�O�kؤts>K�ѣOl��7�&��W�)�d�b�`Q�5W��j�@�RȫVq���B6�Wڨ3&p\�����l��2bi?�Ѱ֥ƝX�&/����;�Uߕ�h1K�}<��.X��;Ƹؚ�;���B�"�p��
��v�e��+�ΗrN"_3~Nx���� ��C��c+Z�I⍞%�"Ue4Тps �JQ�:Jp�Ɏ��LC�a�XzO����Zzy�@cddH��}��<�L`y��l�N:·Q��!�%���H7�Ŭ�D�� �h"�O�ڵ�����;oqn^���ӄ}�	(�fD`��Gy�{�C��V��\�tp���Gs^�H#!�*ᰟ���:���<� q|�=���O}ꒋ�ȕ<S	l�ٵ5::�T
XB����������+ \�E�?�HsRr���>��?������/�]vY'4"`$��BP��&J����s'I�s�=e͕��P* ~]8���i�ƍ7��oqo��Q��Ui��(Gֿ[4*>Mzx]��x�����(OWN��W�N������s!��z�����d��7*�Z��
����=�w��/��D{�+���9�-R��w/Y:���Xj����w��Y��R�%s�Lu,=c�_�hj�����4�I$=��]��ys!o��͋��UҪ��2qm�/�mQ�:��~mS�$�N��L���6«����J6�d�n��^:�x����.��d)����h��3���U�v��@��~�ӟ�٦ے6g��ܩ`(����e�}��O>�$AN����c!��e�"����޳�k�������8H�ks?Ĵ)W����GZ���vb�tؒ�8B��"���_��-�Iæ5�t|��������	Ͼ���s�?OW	�NO�3`/C�-=��]��$����J,��F����W%u�+B���<���֔�	"^�d��vU�ZnC:��i <�{��9|�0q�<��b)
�b��O�������MV{�	a�OBp�#����,{&�JK��-���nE���������n��c�����6>4 kU���^y�0[�l�-#a��(��6�$Ul߾�-oy�9�G#�|q��#[=�1�Y�/,�~"��?q�Y��F�� 6���o�+�������x(+I�үܥ��Q80�99�\
v��X?Pk����$����.��c,�����ш�`�j<C.4@��X�~���$*èj��J����,�W����^�����5F�.
<$�HxP�d��噮l����
�����O��SY�e�w�a8�&8[
�FG�Y��o�)Lp�û(JӚ"��>p�W�[&cت��!J��nBZ�����w\y����}B��R�Ƒ�\I�%<��:���G��P�#�Ҍ�T��Hx���[�^{��	}+I���Tb~�1=��c;w���[�8��L�:plH#�[�r��/�~x�Yg�Ԁq"sĀ�Y�h�?���>��w�3	�`�Y���`c �9�4M�4���'�ŖQ×j�
6�n~�]w�G���P�჈�*�f)�_��W��q���ȓ��<��Ϟ����;�]��p=98&JB��?-�W�	�1�-7D)m
j[���*F�Ņ��p�7)�Ko}�g\�[��*�'��pM'!v��GEV�:6�Tk���#~��ԏ����������rbz3א퍵�f���\zPp�B�Y:l�P{��.F�/��뙧�$�����%�X�q�DNb��֝v�Ԍ�rNY�L-L���d����������1�Ϻ�XgEch�>80�@��USC�q��V;��IZX��������TS�f�j�
�d���\X��#L^c���>�./3�V�FjjXiMiM�;x���Kb���w�꒩ ����{���7LaA����y��j��M�� ����q&8!u�`�J(�1z�Hi�������ť�E�#�J&B�b�Y�^iJ[� �F�*�.���86�iuY�xr�ӣ�v��q��W���~�P1��+)��W��������k���w��_�A��R���}>�я�~��33G�LS{��i q�����o8�����?'dN�q��G��4��ꪫ�Qr�E;22d-z�p^�J��!<~�9�|�#A�UDq�.�*`_BZ�3�I����fI\�� D^�D��|���ymq�uӻn9c�fT-�(f���g�~
?`#HG!ILkN;EO[gpC�h6�lab|�D�v�=M���/�x�ڵ,�R�_lB��Rᙿ�[������ɣ�]��j�����V`�BS�����D₾��o�.N�DI8�k*.��ވɾ���}Ml�l������H�Ǿ�벿2���@�\s�H	�;m�m�)ߵ�4���H����3E��l�[XrY���ht�9��h�}:��c�gX=�DE^^}��7ɗ��;m��a�-�:��4�F���OzYs��!�Q�F�	D[��ġN�ۧ�"��Þ2�lRR��Cj�o�Y�|����T ��UR~#���j*6�������q6�ǡ��KP	�P�9 ���S��s�=���o|�	���|��`.��\"�k#9r��i�g	EB���)�U���oz�K/�D���/,B:���.À�Ę��Y���4"�4��w.�2��Z�͔`;�%~g�R3�aF����$��j�
%M�!k��0�#��^>�b$fP��ƃ>�ļC�����n�?w�F6ՑQ؂�I��L_Ab�o}+����7�R�� "�hH�I3�;H%���)	m��y�E}�C��=:�6S�-W鑚�uDj(��w~�wn��f� 1�JHlm�S;4C���G��N̝f
%nf�
q�������'m��b�t��T�t�S�����[���]�/=�7/!~i��	��@3˞Ye����9��.2��O�|I�c�j�OBa8ܧ4�ۺ�|�OG�*>��֩�+]�d���L��3�S���鮠tm���d�W{���0�Hg���P���78@��iv��Ƌv!k�n30448��wo;&�D�[*��d�r����E�z�6V�W덑��3��p��U�%�$]����Rfڝ�(���o%J62���-��u�����"
�L���3'\�d9b�t�q��c�2|Z����JTx�������7�t�u�]�(�C�aEmvfV�w����{����_�����%�-��Hgt$H1�+�&P�i0����?���~����Z	[9�-w�j-�7$g���j%%������K��#����Iw��������^oC+ Z�_��?�7����/c����4΄#��:$�y�s���v1{l>w�X�m�;�c����|���"��\� d[B������_p����TC���A��Z��&�.Z���>�����!.nO�W�L,ኜӑ�4,o�=�a���J�c݈���s�NZ���jf���.I̐K�g�:i��0�#�<F��b�@"�RW����J|��nD	0�٨�,���z��	��@a|�?M ��4����{��ONp*�[�\�! ��!ĳb�8�r����b�!�}R�S� �t�ZD_�T �P�}�*�� ��flO0B������'(���U�����M�.��TE���<h��!�gT�9���>uӜ�f�L*�9����DaL�F��޸��MNʚO�}�==V�b�O�>���4A�[�T]�N5�2r!���/�RRl�x�,��#J??m
�!�%�^�C>)�i��kR��;�9DL�?̅oI{��W^���Y����������pJ�DE��G}��K.��м��pĳ� P�}{�Y������7�x�5kh�袛�Na0sk�Ə~�����~�ȏ�5ZM��a�F�Xrh�������|��G�-֍�c/ ��Ko�c��������v��"�PM��{�g~���}�c۴iS'�Y�:'��KF	�^�����I�X����B�yA�-g�9�"���ڵ�K_�����6ҁ�(�e�p�#T�\�|衇�7�p��
���V�-��J�$��ӟ>v�y�]~��P�uv0���� r�e|��i0NR�s�da ��]o�>]66ب�S$*�=�vK�zx�Ӆ'�-*�go>���>n��0�$2&b����*�W[6h�nB�˦�i��3��۷m۶={��M�

���D��H-�>�r~�WM��2�*���*g''��p�_��ڱcSe%�؁��A��F�^Y5�&�������n�:�򴝻��=}�k�L�Z���\���nh#Y|Y��7�;C b�:���|>%��4K���^Y��Z�K	�g9���x���hڤ��ԲaAb������2Հ�(7ԜC7�Dӑm@F���)PE(;#�����o�׿�.g���� �;v�{����}��ĕ�̶rHY��/����c�!匸X��*�s �/	�j�&92?زy+�"7G'ͦ�)�&�I�js�X��qRn���.eJ @�e�8�I�Ih������a���n�z�%���^l/�)8��S��9R�2�,��@��{���ܴ����!u��*9�����I�7o_��F��$h�z-d����IZ9��
t��k����2A�B��&_t�Ex�VU�W�'�$�۪�.׍j�p�:r���}�{-�-A��v�����1:<2<8���}/�����޽v5��U�/D.��MBF�����6�eW����}����'D� [�����2L��H�"�,��j�Fs�j����r�2����uúP�;X����D�u�U���b4)��)��i����N?����c�f^|�E�RT�s�l=���v�.hu��.rT�`���+V��W۷������\z�Y[Υ�}��WYhIO�4�|����QE�����Nܯ@���\5M�n$��dOs��KV�G �ұ�Qh���?��sW��٥��S��b����d�P�'!\�������\���wUx�����SӋ�^ǻ�7}��1r������Di��-C�5nf�U~|� Q>���(b�h��a��
�2�5��ѕ���g�:{��D�.�P�I��PRk&ʊ����&L'/:�ꇲא������y�b���{�����,����L��s���_���F���3*��&�J y��/|�������pϪy۫5c"�0�z�j�I_���n��[n������"����CZɯ|�+4���ۿ���u��R��İ�(6� M�����O/��R'f�x5�A�������z��	c�PV��0G�9h$tF~��ô&�sW�]�DW+Ș���_�j�޽4�6 q)	�lT$��5Nsy���醄����[��^��p6���y���n�8�"'�Y�7�OJ4$ 1_����A�� �A��S��u鱵���K�,;�+��b����B�a�y����z���C
�R�\=�4_:V_|1��/~��\:1����O?�j��fbb�����,[���"��W�(��]wb|ݵ犵���y3�N}��X���ܱk���e1Ш��i@F�l~媱᣶e���9D��s��,�YQ-:��m�Z؄�J���;=jÜa�/;�16jR"*�[��.Av���,��W)%�1	�֝�Z�d��a��"ψ���,��P�
^���i���U�+!<�8﷾�-�ozӛ2���x#��!:�u�]`�h�|����$-g�"F��Ց�I��Ç�"���lc�r>s��9�a�kǎͭXQ!)�fՄ�Yc�B0L���>0@�"λ�~����&��Ɖ�X	E��Ej�����Ƥb�H|G�)�������Ƈ�9���%j��᤿�N[�l�Q!��o��<�R����e�)�TOb�(��	�j��C� ZU�k��e�]fC�Yz�N��A�Ҳ�����_N��D<��w��hH2B�U���޽�3��� �c��������4M�I$i���j�_�V�B�ԭM�d|��׾�O��?���_z�%Z��"f%�/�U��8���_�����I�s���ҕ����2���ŇT���) >P:jٓv��ꢢ����G���������ė�H3�n��LB�v�:(/$�ӆ.4����TeD�$��V^Ĉ��]���3	�')�����6!(������4G?�ԫ5�!�9�� ��RL�$�
L��Ѻjժ�*�=�_�rëG��|GS'�g��\E���!h*H��T�Տͩ�9X�臍����d��e��Y�U�X��eJ{Kp�VŻ#�ew4��.܉q�	^z�e���W|]J�yU��V�	J&[Hy6��$�I�?�����#��G�
��������h��w�Bb��#�I��`:��-�;Ｓ>��A����&��b�����7�(	j��2�T�n=><LH��������Щ:�ڱ�ӕI9�l_��W�'�\�`1A!-C�?�%z:)4SXH���`4i�Duk�	��>���"\�� �g�(h��_���rC0k�j%�i�O=��vH�N���0�b��x��g15�6JTU>;;�$<ڈ-��C��E&�	k�VӋN�w�/H�f��K�Pe���в��,�1=9��:���R����9q�+�����7�ˢG�,�GE�`껦�~��Yo>v����j���	{,�!��7�񍷼�&�Ͳ�3Ӥ��F��n"q;��u��3B�N�O�N(�������a���L�!��~�裏��m�Ѐ����^�axD�ڍ�M|{��96��"�Ʋ�l;/O�eC��c+�'قa��r����J��ۻ��=kC+��d}�ThW��pk¡��w���0�/
L�;����p��Y��*�&�YגCRH
�nY���x��n�	^����:��gp��\�|⼰���MI��{"
�wIo$_�*ɪ������ر������	Y{*d2��Q ������3��`�j�m�̑���=2u�P�ȳ��B�ϋΧ��NGF���c:a
����^J�*>FbDg��	��Ͼ��B�1�y����4n��Ƴ�:�H��3NiK�6���(=���lܸ�΀���-��7Q�1�9����'�:������;�x��g?�e���k;�&-lʛb
_x�%e�����?����_O�-��#�݅F�l_���9r�W��A���[pЩ�I��S�<��o�ρ:��i��J���WX�~Ʊ�H,���sσ>H2,��Jz�"��J�}�o��op5��Q�k~�r�ws]v��{I��F|�z" �4ޤ�h���F+C��g]���և6G�g��p���l飤Y�/=�ʦ�n>�❽?b[v��&�ԕ�;$�n���?��?�r�&"��ɣ�����e���9�F&BB>0	�Tb�H>�SRH���t
6�[��~�h�(�nu�СR��iC'V�9c�fR=�w��ب����N�*C6��%%d�)�SU�њ�f�f^��g��<mQC\kX��o�����������F�P%K�Ih^)�f�ې��MsP`��c]2�Iod^��}SúĐ�xX�����b���MW�IE��E�j�bVd�.,���Y�ַ�E��n�:_��C�}�u�ԲTKn_���	��"L� �2o�a���y�������^x!�zB@4}�87�a*�L!e���.a�|��b/��b{�%H- r���?�O���U�'�=��s$l�b�z�\2���������Қ�r�-���sڟ���,P���M����ѳ�g�����/�@�����Ozbb�nnCy?@E؝���{���;n��V((��X78	@�P���鍊n�ű	G:3�	.�,�E��$�H����*���HbF���H���Tk��;[`���%I?��k6l؀�C(D�Ӝ"d�PF�-;�5��\�	(��Ԝ2k=\�Q��"6���+��G��0��!3}�4%�����w||Ex�~z-��$�������I�"xD���oV�`���`Ӎ�ے�#AHpj�Ν$���/���.��гH�J����X6tQ�\��)�k�;⮽GN�	�M�M�.ٸ~W�����o"��%û��fn�ޣ�6ҩ8�f�rq�5�b� ��^�qe��4�N�t�ԙc�Mk���t���4���դ��,��4���E2�����5�^�K?�Y�R��܆'_1�θ�r�*oU��a%!�%�>yx�w֩Q,�X)���ǉŠ�f�4(^�SW�&���G?Jx��,t��� T�[h.~�_���k����pb�8A<�T�&m"�X���ng��q��}Y��J£hͅ��r�B�=~���,|��o�|���~ק+�t~a�tyE��J�K��(���x�{｟����[ba0�"��5��o�w׎���׾�����ҋ��X�2z�i�$Zqǎ���?CmժUt%��bV����铻p]�i�&s֕D{�4�^z�%���Ϧ�/�#MwF]L��-�ﾇz�p��ohԐ�RI*Pt�83'q��qb���.��"b����[y�ng��i:u��D C���8缭�wH7(%A�/�lA~�!u�Eo����,,p!��v�)�d&�`O � ��}�{	liH��cCy�.H]ɍSk�z~�PY���셆<� �㤫Č+~N��!���*���%"��\����0;��l�0�@?��OI��&p�u�ц��ӱ��X�ɒn4}H���/s|m�C8�'���z��\�q�i�]z��;^�Qj0[����-����7ϕ��a�B���5��pv�����qYi��c�E�@�Ni�8˶c�"��Q��L?�z�/�v���J�:x����-;Y5[���)�Z߆��1b@s���e�9E|ݽ��yJt��1N�;��F�Zc���.Z�z�]u�UD"��4¯a�H�~I����S��]Lz�>���håi��L^���	ui��$3p9v;���&M��̿����>��3��M@c(�¿��IU *"�!ݓ����V�7���ox���*D�&���$��O|�	����g�g4*�0���D��`�&�D���&�C� 
��r��C���<��4�?��?��V�����	��i��D%ɱy�f-��z�!0����|�;��������Pt_Q�!������g�����  q��&�S�%�9=��������˯�����`{+\���"E}��_%���뮗"�\t���S� 
1�x�C������tS�{���*=�'˘��k�{���Aw
�`},�kCp����?�<bǴ�����aA�,d�.�B������<Ņ&������k�hR84�݉=�d�mۈ�	�Ӫn��T�+ͫ�Yu�����~J�W6�[�ؙ;:75���t���D������T��>x�@��tq�h��X�D��VS�����<K	X7Z��C	q�	����S�Ă�6k�V����,��Kn��m���een;��V�ºTҾ5e���B�s�e�kD[�p��0��bi5WfĎH�[W�p4�݉>i%oؿ��T�^���5��0Z��[�XH*�U@?x�0��[��\�a^S��W6��<��L�Xl�||���W]�%/�pO&�D��C9�RSht$S)1�5�\�bl���[�����j!�Ɲ|�����d�؜'�}���&��0&@����F�]p��4�L�w�|+{���H�^J��t%�t4�V1�O~򓧟~��i,���0�H�v�nxɃ�q�ԧ�� z�n�t�N�2H�7���k�F����|�iY	��akz�;�I��T~�@�WZ7ԲZ�VA%�Ź��ם~� �9ߴ�V�vy�r�gb�a�9���p�uW����#�j�U�Z�I�b�,ll
=R�H�~�����+K����ޕ��&�H�.�����R��I�����D#cX�mT��Il�}NEAb�C�0-���g|�Ch-%���^�� �q�w3���7�>�~�JeU����L�Dk}�p�8n�j����O���^�0o����chXN2��D�[��ޓ۾��͛�ؽ{��&�f�M[�H�����ʰIb5+5��FhUP���q!Ԛ�e�>��M##Ck&V�5SG��޳��o;�L��\O�!'Z�g�$�iY���ZX���_{vXMi�ʕ$%ff���N3��FL����vڍ�A��`�k`u����9�����=9>�0�h
�a�RÌ	Y�4~ٶ2p�D͚ GE�z�]U"~�ǚ��9!���Z�o�r�R��ڨm:��䧾BK�mWꬖ!� g�=~!2����@�Uw�r������iL��/�ھ�0��}O�ȕ�����u)Z'|k���X`<��@t� e���(f�������i��5t�ہJO�s,\^U�JKe��V}���+�Y�� �Y9u�r���+�bt1\�X��hX��#F����r'�kƙ��t�cqN�B>��7ߜ�U�FJ@�@�Ps�|����?����aT�E�8,fJ����_�J'�+H*�'�+����Ԑ�$d�Z��VC�!��$ǖ-[�j��2�Z+��X�O�ICj��8`lT��({Km�^w婿�[X�8�od�L���y(��v|%M�Ȇd�@�� 6FH�N�V�MUs���cǎ��C]��N�H���BKh�Ы�s����Ms�|��3��������@�648��5��U+V����թ�h�[5����<	~�j��S
AK+ɐN�bl��R��$x�1����:	*��$��	�Jl�^o����à;���'_F�e:)%��,fmC�i,3�)���(���5S	����j��7�����w��Tp%)z%��d�,���(�6��Ui(a��J�]��Ŝ#:���ڑ\Щ�4�� o�]X���$�~����(x܅�j�Z��m��¼��*	��T&xPZ:�0$��p-��&I 3`®p��:�«����4w�����q#CK�K7��*�.d][�!@J�"�7D�%IG�\���s�	̡�#V�v����,�C�0�]�z�oT/V	K74�M�6�-̣6L��X�"t#���݀���i9��8�G\p�@�$�O�g!�[F
F>��i輁 �(6ز�P,A��;����p�k���K�1}g�{M��Y�8vl��H7F��۷��O;�9bc�P��a�A�;�N�Ğk�2w��y�p>|�ݻ��)R�JRG�-��v|�6�ˋHVql�F���R<�TK"ۼ �)Y�'����4D,����9�l�h�@�N�ኖ
�_��D}5u���wc��!Y��fV�~��2a�m��5�]nGOf����\/�?��}x���L�,C�'k9��i$oC���r��!�9��m�����>�$&���4$觾�dT�8D�
`�' ��c�-X��M�C�z�����Z�!�,*{\��bZmÆ'��eo�&�D�2��-��OC4Hb���q���;^����O�N.���� tp�,�W2"��W��/���V�yQn�d��A�dǩP�H�(-�,���ЦRK+:������P[e�t��#�;��]��Ne�EH��՚F�@�R<dC���,�CB������֒��WB��$�(C3
Zp���w��w��~X�ҒC�gϞ^x��/���&)���ϣU.�K׬Y311q�W�������P:���([�os���ߗ^z隷]M�I7$��:|h�`��γ�>�X%]Ϲl>����Q�+�������:U
�"-��FV�y�@�^�޽D+��AE�4�WuЄ�D*֗�v(�B�[�����e="�"�T��8�p�cJx�����knqa0��n
=�M��mo
�;Y<u��M��p��؊ݟ����F����(-�*���)��c���E���V��q��T�fV��R���Ÿ�ej��Xv���SJi{`H)�
���t��fl32U�lj�o�{�a��6ҵ�x�+�uC7� OH�ᕅ�PX��C��?��[F��X�H!�J(��v�Vӛ#�,�@X�]��Jh+����6�� �Rs��+J!_����Q-�
VA�Z��f
��ӌ��+f4��+C�&�V�܏��
���5�Q��6��WH���xOh��+mg&���ѷ��V��ח�ҷ�D+��;:$���%�i7=�f�I���h,�v��sk�#y�L7	�c�\H�7>�����z]|R	��ax!���XE<' d�|ߟGy�ˮM���[���Op9��A�g�Zu.��9�D��{&�N�\�RDTg�g�y�k_:}���^{�.syGbo�xz�+���G�z��یV����.�
k�^<�4�ϧ�%	�(uzn
���4N�g��d�Cj�8ˡv�a�;��8h�Nb?:�\q-�:�w��=��	X�镮K���;j{��I_J7B.1�Ǧ���1�Tz|/"�<J��D=�P��<�)��XL���D�?�����xl��auqFO������-Yj��ŏ���=f
��P�ޅ~�6r�➈��}4�'PC\Ú8���?�, �I�1Nn�ip�O���(�֢"}�U���-���,ɫ�����։�RqE��90���ƀ�kJ)�UWi/X�q"��˨"Rj�� �i]C\�u։cl(��`��0"%:�V2�J`�������CaR��bY�xyT��!a�uF�<K��������x6м��{�n��3�j˖-�7o޷o���k��&N��l�����w�̀�Pca髽{����?��'?I̚��ȅ�F�6�XҔ� �Q��F��� �+��b�V����9|mC|�	�$�f�N;6XJ3o���zq�+���<���W�)A어�#��.�J1���\�1-��w�"�����32���Zv��uG�r����*"�ˁk=r��Ų�9���	�x���Jm����E����:�qh���I��J��!ltp>(�Ɓ���O=/�B��{rFkw��FU*vv$F�����f�WpFZ�O���� �j�R�cp�.�n'�6�o���(2�ݚj�Z�;Q��D�Z&F��������u��{K7+/5��eٕ.��n��
����D�j^�M�$�U>tUIGG1���s3k�%_Ĥ�$�^�|�]�1 ��i�i�^�)��t����) lrV+�K���b�2��`���\P�HD�º�0��(�q���[VF�Z�X�集4]�L)ծ��`��݈x�\��pׇ�^h�UЭ�B�sd>�Q��TO[}.��a*H���������掯�8_"���*uDO~�_$�N���PFnU�,m۶��~׻����ڭ6x}����l��?����C�	�q����Eo��_�3�QD���j/���+�K%�t���R!n�0���!�D	$>/�N2�R>Eu�)oj��A�u�5���aE0�����ǔO�#/�8}w�O|�Y���'��cu��mr�$ -��8��x�w(���\���Jh]Ȍä꯫2*���N�Z3�Q;j���;��J��b���u�>8�F47bmI_�8u�@E�{���[�3�^5��D�s-@�~��
s�Tԃ�6:b�ɼ����YH�fR`\�͔�� E��J^c��*	v�T�g�y�U����##G��#2��l��+2Y��)(T�z�m�Q-a��,X4�xnBoo�R�.@Χ7�������=P-B9Y+ T ���!�� ��NBo�"�	�����P�\^W��O���!�'�����Y�)f�x����H����������nݺ�������h���"W� �����'!�SSS��w��y�m����,�b>t���Ç�������+�C�+�؋�Zr���s����Zпsx$�lt�x^pM��t�f��8vt��ndh�1��ywi�V':��eH3'�*_l��q�z"�o��LT+�y�� XZ�+}�>.:�R�A�Q��*��_1�Ů�!�-f��F='j0��`�ŉ��#�4�=3���B0�C	�Zl�	d#�����-�;��˸�c3lt��\8�HT.��V&E�X�lL�����&s,ƃ�+\
�J��/lY0Y�ݍ~!����'K�:�vk�x�B(ՆH�j"���`�1j���!TF[��hIm�'��J4$N�I�Z(}�N��j�݌n1�.�LJ�_�C`����	���o�;��Ā�u�M*���Z`�LЅ2��+�*#E 
�h#TC�4&	��RbȌ����5tO��4i���w�#Y( �~i1v�#���
�1�Y���gA=���:ؗ����JJ�iwMLz�#����eeэ�2L��$�y�{�������E�q�F���#߷o�Wbk+�WB�+6@���H)�����{�ݴa=�k�*�޽��HKۉj����q��,8����/#�P���N	���nP'Q�qzz���}�E�
��&^D��� R��}84 �b)��y�RMCE:�$����͋�c)�=ޛ��|�w�I�yYv=N�z�!�̑���D��Է���k�K�TIh@'��t!��F��}l�C[Z���T����+7ȫ�8b�Ĭ����PJ;Ƥ�/p[���i�����$$L*�J%�����68�T��C�!q#�n`=: �v�qpCxb�P�-��%[�(���Dqxe�Tz{�M��@�P,�ڈ\o[?
�->Ȟ�p�(i3�A�+�b�q�ƠΟ�&<C�Q�x��N���\aeh��)b!�z�Jꊩu��&����c"��m��2r�����*�%-�%Y��3�k�[���Fu�=��L^tBÇ�8p��0'�0#b���>�C<��ON-��y�X�>4��S�h�=T�%�L�
��MGZ��
bGJ�M{��i�����C��v�ux�yF� ��'���������.�RZ��m��	wg�7�^���Y3q�F�=Q"����Է��s�����m[/Q�/&n}/�D�y c�`�Q^&T��������Q�IwAWE /@7�L�H�
a�a�Q�c����IJ.��T��#e$�o��6b�]�-�D��]�� TT�<x��2�/_W0�Q, `��=�ؐ�hBLs�J"m�Т���p����q+#L�rqq�����5��0�+�j։��)[W=R5�<�mBL�nJ��.���QK�Bo�]�.���a:�n��O�E��Y�p��>��eq���to�O���8W��
�L�ݝ��bX��S�8dR���G�P�g~�k�?˲��7J��zBUs�AS�<�+KD�����~��a�d�^�1肅��tz����P��ө�_� 	lN*%q��~t^��r\��v�<���b�n2M�2�aL��>J��R�"i�OE"Ǉ�įe�i��S��YN��r)M�Ē�&��5���y��B���>�f�5'}������,U�
����c�{p�,dU �$Q��"��)3�z��FL��A1�KBk.e������P�*V� u�j�*�xa���Рߪ�ǯM�%mC̖�n���R��G�t��8ƍ�.�;�D�j��pu��2nB�܈j!V�D �}gDm}}��z�ep{����BeR̵c�K�.��5KN��l����?e��[u�[A�*�.�|���̼��k�TBU�}�T�(B�k�>�(�EXOH�������2���rB��!��:��F�9l|l����*L"��ϭ]��F0PaMa�0�ۍ!���(w�+J)@S��#��i��P�e�Mt�(R����E7 u�銼S&l��L~C�ѯ��s�xz�82�?����/OpEy%��	�gM�0��E�Y�Jb^�t�4T��X]����܍�(	A�Qd�O�����4M����Q�m)�DD"�xtR�� � ,��=�2���0h�u��mUM�+��:A�Vñ��D�>�Tؐ:�\����®%�_A��]�|~a�ϝy��'��/ HU��^j"X�R��N�Ԁ6	~��]�p�Ә^�c��h]���9�Ѫ�l(��Ɩ�$8�:Q���Le�IXL�1��������n�T��!	!&�fe��P����G
�F����1����"���K���K�)_�>g��LǓ����Ⱥ; -�k�+{2��TbI��j�l���c���<n	���)��B�K���^��I>:�b��{��-6;;�F4���k48��X�v�A����1��]	ԫ����x�CI9��}�<��~h{�2�� 祿:�#�\I�3mL��C�]�/Z�=�&��yQz^��`@�X�&�3ү\H�.�P�Xow�ec�z�f���*UX����e41Xg����]����DWU��6
��=UH�DW��>ܳ��4=�m�vO� +�ng�1�&�E���L�g�*(6�����1.��5QG��fL�%G�\�3@jjU9�%P�B��xu��C(�U�4p.#g�*n9c��VI+f�J����� ����:r��9����}Paj�]vD'��j!j������Zv��0U�<���1<<�����Ê��w�<U:�%�ޓ�{�S��y&��:����N�ZiN���K��⫯�:\��L���X��E��N���a���}7ڋ$@<�F8Q&�4.)�~�cź�"q/A�`�#U1$�]�9�I��r�_���Kﶔ�c��m���9��q�UH���FV��n6�?��Y{��w5��C�Z��W	׿�b��aں�Z#PLRa�Q1���GD�H��}/r��M�z�C2����IlOӔk���԰��{�n�O�ڤ�(�&[g=F[FJ`���]h?��n�g��	T�d�����q�<HY9�\P^��|�6Ī�OW���95�ȋƆpF@f�'�>�`SmB��<ʯq��b"I�ԥ��Co� �*�u�u1غx��1w�1|���)1��JDk���Q��)�k��6j���>�6T蝙�A��$�cl��8�k���ϧ7۷�ܵk�<�������/��g�i�$����!�����5����o��{z�t@�.J���_�b�m���_c#������"�u�J��g&����3��q�*���{~ ��r�<�c:��zyZ�������Y^D�S��K�y�W�~(e��%��iuQכ������a;4��u=�z��s�iȆШ2=�`�Yh��^�؜���D���*-l��ۄ��Y�c��n���+��B�\�����kC �ZK�Q�V���j����ֱ}\@��LE@ ����c�	f{%���E�ʐ��d?��6�O�^�(�
|���j`R(&��I��*h��R�_4��y�fJ�u!r�_��l⮈=�=��@t���Z���鋊�	�z��ڄC�e��z}J؈!��R�cGW�~��Ui�I�z͚5��8��k����c�&������u�Y�ׯ��h;���w���?>P�^s�5��}�����j���"r�.��^6�E�U�B����_�坼��V�ڠ[�ZѨ��C4�vs��щU������+���^��y��F�,��zh��ZlUO*5&�$-���ש�ZWk�1y�7��a.O�V��xU�rv,	��ld2���c�z�.c0b�M��M���B�e��؇�lѓiW	MtMz_�80\�:��VSo�H"ϸ�jAW�����]�F9;Z��^���p�؅��Ct��:$s�����*i��Z����sq>�Tk<���f-�I�2���k���Riyx�e⃑S���+��(}����c<+Q��a���+��̆jA�D`*E�=����4I��ҵ��Х0,���sGn����W�H�H�E��1�X]b�y�������l�srd��kwڭv\��9g	J��&�>Di��X]��(-{�Z�J�0���(��w���Ӥ>O����@o!y���WZ�N���"s��EҐp�
ت�1�i���$�6b���nŜT����D�5`�y����1J#;��V�7�b�5�%I7V�Ke����48P�r����8��O��k�������D8]�MLL��-���|��yzz�h��f�q�3��F���>o��'d+8��IV�]�a�Z��?�o���o\c�F���,�s���wwݺu�O[M����g��%��&������X4��C���	,#	��I4�a��2X�,��4�
���1��О����L��Z9k!��#�F�b$*R暼�Y.|ʊ�_pNA��)�Dm7c�����
��jX��A��k)xW���.���4D����TLD�G����A�:/f�i�'�3>��ˉB��1uxY��m$7ĈYY�]��*K���Y��i(�@xL3�֝��MeĨy��I������jM�����g��(Ӭ���>H���n(� 
i�g$����B�&Ž��H6���G⦡ox�%��vk�+:6����$��u����ꘄԬ_m@T5U|nK�����z�p�k�2ʸv[���!�3�b���:��q����Sl�v>��D�w��+�P��~��1�72>�x���@�O z����5kV�^�%�0�����/�L�s�A+��cs(��8��g�I}���pd�`Ah}b�8�j��}��e6- ��r�i�M9*]�8@�D�# �b?�S�7�$\%)�i٪�,	��F��/̷�g�#��S�d�������k�m�v�5��=ߨ��e5"ʼ�5|~+��h��ڄ�U�Ɣ�r�u^�A*�?%�6t����+EO&h�}�.Q�O�(�ŁĴ����$�Iⶑ�:�H���a���k���Et���%I�;x�BC9���Z�*[ɥ#��>xDt�n�t.Hq��}\�֩q,6�d�J;㞅� I�h%������"'-�=�Ϣ��&b4�	0��G/Ӆ������B3�x�\����bv��"ʨ�a���&�J�n���x�	G4/�X�/B�v��Mt* 9�o��\Y7]�������z.t�b�U���$r<�G���A��\�T3�b��w����=�\Jc��b�#Q�B������L𷡒;j�p�E�	LW��^96JLx���t֮�⊍7n=�K>�vJ�uϞ=۶m;p`����OL��r��~FV����京$=�xt���7�|��I�F��w�O~�f�93s��''3D���|A��ˑ��bNT?�H|�QW,�$t��Ѹ�&''W�X�ܠt�[��os�H��X�ڒ,����1q�5Ľ�e�g.�p�'��^&�m��v9x�R�0A��Rf�~�=w�+�j�S�3�<H0Q8��@�2*���վ$V�h�R�>N�Dw��J�dV��_��r���"�L��a�v�Q<lJ��HO!SeU����rNϪ.2�v�-�Qɘ���`�1���{+�e`������5Kd�y��&����5K3`&BFD���T��(�֔e�M>L~��ֆ�jY�Q4��'�� �A��V����YF�~��B�vl4O�����CnWJ�Ȕ_���t_��>o����Lz�u;���n��MK�H��.��7��M�~���w^j�S��.��n��+�<�����><	X�󒰵J�'$F����3���>���������Q���U����}��ĵ��-�s�H
V;���H}��~f���ʢ�孊q#���l7�㱱���t`Zy�b���+uֹ:9��k������6b��Z�X���#1�V��	<�l�,m�T���k�ʉ5d�v�j+���r��*�'��D�d�F�J$4���ZO�=��b	Y�Y/��r��#0�Pw-	\�4�^�GPMMe���t�
����#��)i�H"1R�"�/���D�	aP�Q�g��j�?�AiB��Е7x��}�=0�0+R\�O*|'I(`d�D�إQ_1�i��.}����*U�]Wcq�]7�2E����� o[N���&�t�'�%]�������p�H���FwAb%!{ȅ��j3��T5����&z�+��t���N@H�G��qYH����Je�KO�.$��AZ;,>1�PxdBXKR�U���v�e<�U}T*,����2��;�ep5-���舑f9Ozz�ٷ\u�>���k�����^" <33C�{ӆ���֛n�}�����.Ոױ')ʹ��cǪ����=�]��4�z%#��;�8�ׯ?���}��5���֨$4G�l�1AOeS{��6��lN��<�`"�ɛD�lvvv��~vr��k�L\!�~ʎ�iUj	�� ԃ2(�@̌�-S��Z�^��siw4��G��W�%�Կ�K^�fw�Y����Sz��4�0�#��vBg/�.��Z����S�vPץ	~|P<-�����u1��OU��Q���L�o��0�M�#1 �u��L�g�S�IA}ō�*�n)�x�lT�+���'I�\#֢���Ԩ꧘H�2F��gP���_�}"cl7��F�`����I�VNBN*�d��Q���"Ҋ���Wk	z����䲪h`|�w�jy�u��촕��i�U��q�Unt��L16�?��9Q)V�v��NB�;h�dZ*�m���IC��ƉϦҒ�dJ�F:{1������o��F�cccO<����� LM�����̍��q�[�n%�=��x��w���Άj�}r�uW���o%�}�>���'��œONOO֦�7�~����؊ї^zi�W����"�Gj�#�_V#�O)]6�科�hX��9O�900D�g��Denn��,��ǉ�g5��`e�"Q"�z�������ə���׮�-��Y;7��S�^f����)K�[W��tE)��t��,��_��G����{�k`99ˆT���������mW%����h�QPs����w����$�$e)mc<#�]ς�ְ��r�}�0-�	�s"�4�le:����U�V2(z���< +	����9"��?E��E��w\ܭ\��xM�1�jwV�Q>^	ţ�pܩH�U�-�hz���zܩ԰����B�E��w{��ݣ̢k���n��V�2U����'}��M0������� ?A,f����\@$����m�u�㣄�wE�.����v�����'!�^5�y�u<��:����ق�Ƨ��ަk��ӛ�+V�}�9+W�$��٧����H�vddĖ��@crr�{���+/��믹��=ؖy��\?��H��K��/�馛��������/~��67t��C����x���~����|�����/}� |�6��
0!���x���/�B/}9����|��V�XAB���i]Eb�Z$=jc��1��#u�F����D��FΏ��z�z�%�v�����S��D�*�dn5%ED��qU&�%Hv�Kol�ɱ�}����O\����Y)�'I�r]�pC-���l\�e/�Au��E���`�T��t�X�SV�Wܐ5*�+��0Q�x�������*�O�{��ݠ��cB�f�[C�����������P��O��$��V���;�)|:Y3�`����}ƅ��	�[wP�P��SEW��B�!���GY�.����h��VC%��!�կ`B,|���݆ X��0�du���W%�J���V@�����nj��+��Ζ���]0M�Jֺ�.�����۔�nJ0˞M�6�M��H��r��ظq#�2�T���w�`���J%��d���g�}6}~�������K�����K5�����w�����]���2�.��_����_x�������8pB�j��FF�%�vs*���X�B�i�����A6e��V���\�&gMN�侓�ΎiuЗ�3��*s��cGid��P^9�W�8�2l�q�4�U:Piɵ�\�����Yɣ��\�e����S�P�ī��U>)��J�u��n4���Q��2��,�����/�b:���^�Jރ��(#���P��\�P`>���`+�\R%}�#�h���~XK�k�O#An�$�*�9m��F�2,�1��QkI��Y��yN�^��OD�E�T��.�,��6@�L���b�*\�s-<� p`M��p+l�EA�
�]�y׍^*&�A�UF�S��ږN������N�z�&����{�~mB�r�y�Qm<,'I�	+�T�F5���|�.�v0+ɐb}a;h�rZ�J55E�r�f��~��N��t��P2P�KYhQ�!�hY������' 3������r�-�=|?)0VD��v�ۧZT߷�EB��D�йX���I�լ��׮]wlf���)Bӛ6m���ˎ#A�}>k*��͛����f�u�4PrD^V\�� #�<=�j�ʵ��!xd���ÇO;�4��+W*]���U5q_�<�9E��nC&�����z>;Kb��h���'ְf��m6��u��fpx�iɿ�'�?j�Ϛ�:��^������s��F���	@�0��{������R�gn��P�@\���5���~���ڻ � g�k�VrqK 
%�orli�z��`=���p85��Z `�x&i��h����F��J���Bz����I�E���i�x_]�ed�֓����ON�'>i1��+��ݘ�X����*C�n<������\7�0��o�~������k�zmb�g(��=M�=apA�I��t�Y�������e^Y��LQ�k�͢t�4tqsQu=d�*�)+3A{N���x��ۨ����r���(t�D�	lTf$6��>�d4���MCp��V�	��}&��ZZ�;��D1�{H6H؟xѹ������WH+��v��+pl�n�G�j��c��l��G�y������'i�C�����ƌX�`�ͰC�=��xF�z�~&f=8��l2����!B93��<DϦ+��o�x�>ZZ)�i�&���"W��:��󯼶��������Zb������3|���ˉX�H��V�������s�U.�LȤt	A�"[<���Q6������
�]��DLVU�x�O�r��~�G(K/���F�Y�@�8��MȂM�K��.P!��~*�*�:�"g� ^ݓm�����&҈���,�U����'�H����+�=Q�7h�D���!OBr�JS���2��L
CZI*��IQ�2Ut�I��ΘkZ��Z������hQ�[�����^�)���_�4��;�Ҟ��HV��E�┹D��0,:1�S����\\�Q����*+���%'g"J�I�fR��ӫ�ӈ��I����)�(F���$�45;�h[�;�B���,~�PI��S��F�@%��IӪ�z����雤kW��L�R����e� Xa��e�ԙ��ѣ"w�q�fRl.�����[�jeV�f��Y����ސ���)�";�O0�����&�L�P�a�H5D円X-�t�u��OE�߲e��/���\�7����$$r�r烶�h�Ꝅ_#[_4>$��[��CX�V����5k���Ornnnp��VV��f9j��;���4}�0��'&&� �����R��M%
%�eZ3Ɓ���y�Zse�f�3�Dz��(FYC옊Y!�d�[�\�Y�8=��v?\*���vI��$�Y
塡���y����I����R��`_Xw3�S�#�nu��GLQ�q�Zu�F�L�Qқ��&�tA߷�m��_e��v��u=�(�C�J��M��`[A_�I�2�d��˫�.�%��"�W�o��p��2�!�$)�`���D�ń����c��S��}�˘V��R(�R�#�q�(���e��|���Yi4�nܞ7IE*��cE:�NhF;�](D����.T��&�:�2ʠQI�i�@�T0_�T��\����⥟c̐�O=�Ե�^K��Z3�x�;v����O3⤴`��[����[�6��;v�Qgz�A֭[G�&NؙX"���;W�^={lBb�XK���=m=�w�5�LO۹s�#���i��O��n<��`)Nsz����ܱ��3׮ݰa����5��FjC۶m[�])+����ko.,�f�p7V��c+V�:ғ��h�N�LQ6��<uy�8�(�#�H5�n^=;?8x�>1RVRI�/|xyo)=���-Q$wr!���S�J���Bu�>V��~���A��<���z%��l�cB���K!O<$=0p�QzJ�g��*Q|�v��Q��I.�[�+	�;. No�Y��qe�N�$4+}�c�`W�E{=�ȣ�o�;�L���6QYT뵈*��G��,��ͥ�,�B/:E^����<Q)}8==��[u<j����C5wWn㓌��%�#+�,���j D�ؤ&A�j�z������w�,-�	$����1|׃7V`���a�Ĭ�H! kl���/��kM�n�cY��Z-l��٫gP�0���k�2�ΐU����V��Dz��e���M��2=�k����,f&.��̗8��>{�u�M=p��7�ؽ{w�a�OH���/߼y3=��|�W�����o�v�k��޻Ge��x��?�a�e=k�֩�)*ͪ���斔��Ī��ww�~�y�����B��r�.=F�E�ig�]1���_��$q(�B`�����٦�A�1}^��� �:��pԊHl�,�zMBg��]p�ʲ`:�-"���H|�[]`��Ě�<�x���2>t)�Eзt�(+?�=�ܭg�����x�����yTnT}5.J�0AaT��F��$����$�~���_���q�B�l�ee��A�2Lؠl�a�H�X�w�M��x�5�5)���zk�.ⴣ�M4rY]��t"�4�"�m�\X��`Tw��Σ$u�}�ze�ά�`���M� ����!n�o�w9qN�SNWÑ��3�]1��	���dy�] ��v|�E�1��������VcTU�ou�Ph��$�"0�M<>t��J��<˖�W��`�R�>NI4�OITۚ�L8����"6�淼�>_�v�#G&$�!�F<���?��7��vKHբ4^��!p��O^y�o~˕����yF��'i��c+�+[�'���#�N/TOB�dɗ�R�P�,u�'��e�;nQ�1Ti���`�*����ѩ�6nx�׎��^|��� gy����Xɑڦ���ls�L5��'�#l'A91�t;=?�uYMA�b�*U�L�d�����uY�4+�P��$���N�`j��p�H%G$S`C�!]�!x�?��i�a�tl�µ�D��$F�1/[��c���g�>�Oi�
.	3�G�{��ѐ�V4�G�� 9�_�m��2�#=Fc�5��(+���C'�{��bd靈&�yj��`|�[R����F��V0 B>�(�;D��r$��?6Q T��N��6*i��1��.J�1Ar�.�X����E>	��$Y�Asc�P�B������T̢r]�*��mB�%j�ΖY�`!f�&�
�(�[�*��WII��-�:���	�Km�t)M��& �#��fB�6&�,ԱPʉ�j�I�d#1c(A��1���Q� I����;���_����r�-7n$�e˙<��m۶������˯����$��ğM��ߞW��u��.���5�OK%�r������n��V���~n�{$1Zʸ�[���O]�b̄��*�V~��%�p�ر��6h]8�:}�}�>'�JZ�kÌE�ҳ�ryJ�{a*�y�F�S�a�U�W��TX�>E�T᳔KZ_���>�Ly��M��_��C��/q̦�m���y{�hɪ�~t�sNUݡo��Mw3�"A�ADQ�Q������aVV���[�i�2��Z�y�d9DAF���B#25s3446�@�}��U��>��9�[����n�%�,l�V���?���-
2w��R�$�iY_�4�jh�=*T���� ��(��\����؊�$�5zG�e�}���I��&��W�p�v|h�=f`�t8*dtLaQ����,
�$��=P:u�eJB��-�%��㧷by�%�_(�Ҟb@%�ʫ�y�dR��o�nƫe��� ڢ9�C#���-���Z�@*y�,�����ϕ'�~�JD�^|:Tf�a?�l�Je�u�ԴkDmŦ�����*�4j����P�|�	���ɑ7�T�Q��u�L�0����F��4x�[���%����u��=��C6l8��#�k�j>f뛛�{�z
} �e�W�%B@�Z�q���}��+W�<d�ϰ�hc���7�v��?���9VTC�k:��~JJM��(��k�� J6��nJ[���M&����ut�E3Ӳػcd�k6w�l��Y���h�����jP;X��n"�Tzȍ�|�-�ZO����u�],��u*%�gͳH�t�]I��[/ʽ�Hm=o�lr��Ϩ�$����1E���*!=~����TV�J�����5�d�e^4���vJ�g�1=����)�ۛE�[�;7� �4�ݜV�fd�E�)�&���1��)")k\F�F\�OT-��~o�`����6PU��0c������Ĉ�d���jW�M�-�5��MBZӐ���ug}���1n��S��_��¤��d�������ȥ^��&e\>I�� �=)�}ʊ��(���شb����邞L�5�밷���i5����������[�͌Ma��X�zcM����e��bX�?(72��́����ړ^��,x��-�r"NJ�?�`N�-肋������� ttch��j�EI�-��Mo+�pڍ���Ϧ5ᬍ�A�A��F!0�V��c��Im�h��aA��N$���k�����Eo<	)�§�#%ƞ��D=z4�G(�����a/匍��{k �(Ҩ�1�i=�? F䕦x�$)�Y�%�_�@�@ʧgiݗ���m���Gƻ&��.���i����IHdo�I�����I���yC������V�|��]2��l�̙s���]^@�O������ז��{��v�m[�l9��.��2��z��o������l�ϫ|�9��p{39W*�8t��5+������B)v�A����I#�n���lB�#19Y�T� ��Q�9n*ݜ�6o
s������iS��n9]L�{j�Ny���뿱X�r�	P�t띉Ѷp�>����Ѝ%�Fs�����0�ԛVD�	�e�^QP>Q?!}0g�DG�w�
�
%�������.'�P�N��4�3���Hw?��㢧�_�f4�+���}�Ul߬4�!qrzPˢ��vQ.:�htt�S�}���y�
��Y�%��<1OB�T�U9C�Ry@�^N!1�Q�,�	b�t�j�k'�q�m�)bϞ=�`ێH�������ϖX�D�e��R)GUj��ui�������X�����Ӛ����q��^"�5Ub�,J�J�"5�;��U����6r:��E�+^���=�!���@���sfꮈ�iۧd��^�}|6un]�`�����3s��a�Y;�Vr�ѩ��=+a�q1���6m��7����&�9s�J�;#��<�\dL�Ȓ���3��ώ�bo;Y�pv}���䏏�CcI��dɸh?�\/T����5�g.�ܮ�� ��w�2��r!H8��i���t߾�`m`���5�%CI��w�],2��Z3q�µM�)�|`��PM�"s[L�^�V�uvs,�c��+�=�B/���v<�2p����)��6�˘Z��2����~i6�V4$c{'TZ�M-���ި�Ӏ�lԼ��=�Y�ٻ 
e�K/�`�q��*=g���s�IdD�[������2�hvb|��I�I�I����G�����8�r6���0T��t�X{�Ԭ)]���C�<g�d/���$\�[F�{\�܁�d�_�'\b�q�%�"��4(&�SN��S,x&g�����͠M�.&.n1��j��ܒ��B��RD���Q�Q����*}��0�F>W���bP���Y�
0�h�9�!p���KūbZh"�B�{V��I���RO�A��JEFr���B�r�sJ�� 1 ��| ��^0v
������6]�(��p�CX�*D�EUL �e8�|���gU�"Z�&㜊������Ť4��x.����2�ѶE`ux�ː����F�I�������P�W}Dr�6f$>O��N�T`��ը���Lv��"�\��O�P�V�3_n�af�	�?w���&c%�fM�J�V]����و��0�&�C�%5ݞ�0��՛B8�mq��L"�����0ox\\�UC�D�n�=Ri8(�l�����`�I��M,�8V�O�$�/zcC��S�K�I>:i6�I94�1;�l�:u��Q%@�۰���Ρo?�
G�夡�@"95�BݫӐ'/ɪ���g�V�#�(�/a��,�$��C�		S���%�n���%pE�,�Zr�T�u��I`8k�m�P~�M��|��*�\�.$�Hk�S��e��F!��PI��!4�6��� % �+�UR�Z(���Ϛ)ڶ"�t�Qb���s�,���J����O�!�/w�@O������ܒ�p[���v=t�pDaC��x��Յ!�6�~�Tǧ��6"�$���,f^K�v����_ۮ�v�R|Z��r��93���b��]o�ܹsΌ�E��s�N�u1dؠ��l��9ZdIn�b���i��}m�vs�3/N���1��"�,�n�� ���[uҋc][hޜ6䋱ڡ�^0c΢2hzF	VT14+�N���y�o4��+螣���¥��I8`��l?��*D%D]'&^�X�࿬��]�v4���R>���'�������g���^�S�s�Jyy*�o��-+"��&��/�ռY��op���~����v�e���tP�ΞX*;��Q�%VUD����YHT����;v�h6[t����#f�����)�Z߆r�?m�7"����`f�m��_i�n�0{欆(gy��!�)uGQ!���P���=K>)�x�Lx���V$Gbj�=240�����/z�I�!/EVȺJ=M[�Y�C�"7b^��i���ׅ��f����v��/nذ����A!��w�q@at��-[ԍ����6~������xsB�=u�zd��NN6�}�kr�zVC��xA<)#2_a�T�+$�;8՚�g�uӪ_͔G2�IN_�JF�L$��̚ȭ��k�-et�ں������`��	�9�Z-	�r�2-Y���Y��S�m����z�Y�	5��g~߾����l�1<d�b�!򂂧W]�>ĵ�a �]������N���K�7��S�q?�iW�	��DCr���=�Q��B��n=��w�|�ɋ/���h"��FW�l�:�)�����52e�����N*/�"���q�x��!!����H������뮻��B�Y�|�%�\r�'��ي�Y�U�V=���8TE��E�v�i\p���IIƠ�{����u��;W�\y�g� ���(�#��5Q�c��9�l��
z���Ͽ��[i��x��c�97c(�d��Գ�F���R2A��{�+���K�o�Ve�����$��I��=oE@��y^�^���;;I�0c�̋.�ˁg�%c;�H�$�0�2�)�i�)M)�:ɔ��t!���@
��Ф�vՠ�"c�L)����w��]���~=��w}��_�?.���?��0����|��_~׻��>[��LTv\o���rq������4E��@�@ԥĻ����M�t�z6X��W�'�G,>����"��]���u�U�Q"�%]&7=&����!������X���	����9mm޶m����yf�H=-۾�S�?3�8|˾|�[�F��s��֒���"��M#O��g�����Ȝ�0��^)~C�s���d�����#��&i`R�A��Ļ(xH|���6Ơ��8�HB���*�)8�$�t�į�HU=q�Ҥ6<4�C`�斄�H�?�g�Jy���}� ����/~��j�` �#�}��.��������O<�������Z�b�#*.���gϞdA��=p?~��\љg�y�{N�t����)��g K2	V��L2�[)��^"��Yf���֯_���衇����q�?��?~�;�	��׻	�N4"�����UgXub.�EpD#O;�=[[N������XI�.��I��wh���6�:%�?>��� 5*6n���SO��LV��f�e���;��S5�7��*2�`���J��IUꌣ��Φ#��m����ʗh�x����PG�I�'<&��;y.h)��η@`��4 ���51FϦ2�v��v_��Va�A
���F|=����(9���Q�
CIg_�����U����=ǹ�R��Li�c¦^F!Z4�Bf���wFĒ:� �{��C�i�����)��\�� �`��~կE�F��A�mPh����������ζϛ7o����߂�����92R���VT�(e�t�ɪ��/&X~b{ �%���p�3��F��x1�sO3�v�\׿(���eJ>ݗ�2�(i�O�V�5�R���@������rT�;��x�'�|L�\!�s
�۾}{-����w�}�6mZ�d�gI��(%�����LĽǉP��I����Zm-\K��C�MJ�T�sr �q����Xʺ��o���G�A��"���kW^y��?�y�x�D�R񃉆��6���\Rٙn�':tt��G�NT2F�y�)����'��C��<$kv!˾���Tp�Y���o|�g����B`�8��< ��]�l�QGŚ��5���=�^�c��b�![4�:��e�Z��<��AQ\�!��P��:KEH2^��;�p�1Z�q����>A�\�,��`�H��x.j��~�@�'	��T)���Z=U;Ȩh<�Jl��ۓ(����n*��țnδ��~�V�bܦ��U_���Lu)��4�&�FK�;fҝ48���*�9��ң���㵷�'��<��r޿gll�/�>krx8K���_sxx���$���q6�j`x�:�R1I��P"�+D�&Uc\�W4-�㲲UNd^�-���U�&�@��ۅi���=��f�Lg��Z�F�+u��+v�L�tA����K�	g�C翪<��Vl>-w�{2�J�P��w�8�::�sE=L$`M}HRu3�(��yr��"kQ�S�����y�k����A��.���s�p;d���B�	u�.��"�=X���	D�,�j[i TSU|�7��Mo�_��}r_���7�P�ӵ��o�=ЪDy�M�r&�+�l�g���B��Z���I����W�^=o�|>��C)�W÷U����|��b�K/�DYG�Gx�T{���@@�s�9�mo{�\���>��o~[�Wh}�~�ӟ���^	�T���J��R���E�ԏ��Y�g�ݣ���MV��t�ι���(�yd�7D�Z#^�'W�v|*pXS&!"+8�TsHU�!�h�$�����BA� ��H`+�O�]ب�+���E#�%x�(t:W2`Byg5~� ��4�S���<4:�z�m(�+TC� ^[<L�>!�3?Gw�&�/��@c��YJ$[�X̥���Y��${����6|�@�[���}"���Iͬ�H9�FUD�~J2)HQ�^OY��ʈR��p'�޲�����3}�|���G���M�w��K�ty��1��Ը)�`PT��é��i�KlO�(��5s��@�Q}��[��X��3�/��2e��o뭷��4���'�j8�7  �s�#�A�xGj�̞�S��
���Y�f� @̝;�O���X��\���D�hu��Ty��_y� (�閇gɏ3�p�9I�J^.�]�@��|�
n��K����Q��h�ގ�yFHqd鈉��b�Ǽ���Y���������q�� ��Q�?�N#��R2�=�F^����!0�����b�V;�2�NZ�6��G��4�=�NJ���R�1��ڌ��Pe�5�t�����KI��A��{uݦ�LyZq�G�3��<�c4��*�r���U�0�"����r���-$'ެ�̽��]�7c�47��7��I��|k��yf���9w������8;[{&�d2���0X��lm)��*ж&G�`���zn��dF�'1)��N�Ԗ���9y�Ĕ�2%_�}-$..�ZAa��ٷ0�+u/���F�?���R��:�3U�1H?&�E��J���R�L��Q��D�=��K�sf��Dp�C.�����c��z ԟ��F�[ML�ϙ3�]%�����2����8묳���d>�Iun�%K��f!s��zE��S����&�b׮]�>�l*��Dlh�*{l-�Z9�ԤE��
2�[W��p<Q�9sv���o����p��u��}���n|����z�JjMo7����ib�
_f㲖Jلz[|�F0����q����nbp ����������'��ꪫFF���,��>2�2���x�.j`����5�E��w3H�`cH�rfr�bJ������g	fGO��P�����B0*��<pvRf;]����hL����@I���AG@�v��T�4������/�}/���P?�9	�wسg��ٔ��ݙMeMKqs�#iU�U�3��kvfHa��&V���U��b���� ���k��� ?���2ٻL�Ȯ[�g�rCS3W��r����p����/��J�#�����>�6_4�Gw��=o�!+W��.�"��{�=9�ó��,�`��hS
�x�w���饇�2���H͢tE]�-.]�)�Ok�ٷZ�4D�!U�1
�eN�<5U�&�0/���ZH����X�����
o��r�����O_~��[�nÊ̘1]�j�U�}p'D��O?�._N�w��W��m��&3�nP>�ҕb�aCZ�~�෾�-<��0X�C����^�ͷ�z�!�,:�3X�����ZE�X����"��I�� ��o�F.��������!�Q���\r�h�B���'O8���;�8ꨣ���M��������SO5�i���{��!��t1��jZ��I��������S�aW��Pj��C[I�ٚ�Df���~R�]��'|��4~�m���ˇ�0	CC�1WHc��;�o��o�0��k��FFF8�e��ɑ[�XD]��Q�A��B޲��ޛ�W:%���xu��z�t'��5ӧ܈9��O�A��u6��7��"��Z}��$�D"|����ȴxM���̖�^o�g�n�6�}���.8��PO�w ��ld�! �;�tN��n�:c`��m��3�n4��y.#���'
�~f[�Y8�}L
�RYÆuE.����"/�Z��Ĥ���ݪ:[1�~"��ǜu���ni#EU�M��N��U~3U��"��W�XE��4��U�:q���3�y�3y�s�������+�/���y�7�|�yP� �29��������~
�h_�r������9ƪF&qժ�<y�1,@� �����,[���۷n�^uՕ{���*/E`2��q�G`t̬[�U9A�\�y�7i�7O�{B�1�GO0lT�{�P����c͹zmbԗ��,�ҀP�򥉢-�=���O=�=5I'�v�Z (Ue����ܺ�~p-'T����<�L���u�;ѳ�u1����f=O�� H5c�����gZ�%�K������Ql޼��^pQ��[�z�g���+�h˖-�?~��ĝ𕕟�K���7'[T��u#U(h�/z��/�����&�|HK�i��8c��}��h��%�/��vI�w���t;$��6˟��G^Rt*���&������s)\�3=%�O'P��f@�|'��t����	�a���D�$�:P��YWFpJ�כcN9f�l��pAQn���o���4)�f��ԡ�N���WT9t�����D�nŊ%�{�̙,��C9v���~���ڿ�Qi��'����Y
GE''N;��E�*
#�A���-9G*I	y�Ry�!zs�K5�M�;�iT`1�u���Sg�ՄR�<^��3͖�F�FԈ*��%���@��]p�6nܴi��ȅ	?餓��c͚5w�u��B \��ԥP��ıA�@$Qz9:!h&n���{�\u'����I�L����;��1���-Y�$o�]H�n��?"=��0�ܰaË�'K��^
�>����O9>6c��_|�ENf���MGg��ƛ�f�>�(����ZU�����s�Q9�?��ҏ�{�d+D�M�m�Q�c�U��w�$�i#�W���-�6��$p��[n�ă�$2ѯ����W_�@�f���җ���z衫���:�L�Ӌ/��g>��-�S0~������C��5���>���K�*�Е��g�Ĥi4��Ȭ�;w��]xᅸ�Q#<���$۶mC�1v��_oE|����O3C�US�ZZ���#��f ��l-Ŕ�*q�~�s�-��a���W%#���)�k=�:
2�����	���f�ǵ٘�]B�+��C�'7E~����>��$�3+ű^�`�1����&`�3F�[����t Kf�|(M�h��G�Cvl�Mz���x�\���躆�r��	�ۆi!΄�e$��,}Bjm��e}����pڍ��t�4XR��k��ob�%\�R��$<'�f��b�)�C)�/�|j�W��@.�xE��o^JTE��{봠TYU�fd�J��-}���m��4�l,X�H�����f�h@�a�T�,�0
�3ع���ԽZ��%_s�ͷ���=2[!5��<��s ��۷5��_|������ޱ�=��c���/v��U��?�����}  ϗρ]��٣?r��e4�q�����ܳg�}��w�u?z��0`y�	)tTƣ/��ғ�<�[p^k�hHE`�YRx�-�#ɠF����)E뫤�r 3~Sx�d��sf2�D���ˏ��Y���|��n��]e��,��>��Wֿl���2��3�񕍤�"�1���	�n��j�{�����_�ud]�1u��DS<|� ;P@0'L�M7ݲq�F��F��<^
q�*�ΒP���n������Tn�rŲ�=ڶ��|ph����|�j��/�.�b��%�\���~JRYH���M �U��CsG�,���L*�g3�5�����U�f�����7��W�
���e����Rr��º��q�NI,ۍK����c����ˈ�	�1�͉	l�����ص�����>�YMsܫ�F�	j:����C�/,��r1��$��;��6+�8v��B��v!I�����0T0�JC��~
���7�VW�2���������ƦQ�^�|�$��WFW}�~�,$��d�I<��Wd@���:���:�����K/��M���*�FR��$���x�Y�^��iEȏH��:P��^!�cǓO>y�EQ�@.�Z�j���8�e(ݍ-�W�<�o�mL
��O�׹Qgz\����~��/_n��:��dަF��|	�*����Փ���6y��_Db�F*i�z������-[��ٟ�٘T�Ik7'��VY:�
p���ϣ��֚:_�����~��wԤ�'�U.�ܨ���A�TG�'˖-�SyYaַ��$�?�z���1�?��O�,�����q��B;����v��~(�� ���Y��q����is'}�����O�*Y%D��±������ ������_�K����˶b�I�e��n��������x8,�������]����j���IO�W���&���ξ��	Il̬dBRF�V\����f���ji����Թ���ӹ3�f���㧎��]LN���N�{=;J=�Vgf���ei�m;���j-ϲ��N�v�����^Җ��"�t�u����j#3g���d2�.�Y�g2�|g��#YT�ʺN�v���Q�����cϺj�Jc�a��&�| ��ܒH�lW9T��V���x�g]6�,�wJ%^�.��b`�SjR%�(%m6��+�[��K�q_wq����uG��V�$��_�͉�_��G�������?\��ѻ��ghPp�;�c8@p��w�� 
x��o�!��Έ`-J�ֽ Y��HZy{�� ������˗.�18t���6��A�cj�zZˆfx�6�f덖��~���[n�実܁Ύ��$oB��1._���^��i:����쑙����'*�������(.Y{�9�֚�)} "�CBm5�Z5��3W�;���λg͘)'^�e����6�`I�b���Pc�k��״͢��U�9�L}��8�s��RI���<^�v�H ��+�N�X��*9��;�|��5sgϩ�oy��Pm�ZiH˼��}h��'kh�ўl�<f���C���$3��e�1��_�К�n�i�[oz� b��-
|�M L蚧{�����[�'�x"�9���fs�VM���0�l���髥5'N�y٬��ږ ��B�L<�R\�ِ/�aV2PF�sy�#�o�
t��~����wg�9*��u�o>�G"B�:Jp�)���������#�C����u�3��8�f*����x�xb|�'���s��_��h˧zù��Q��NU��+[��x�C�`���+:��Xِ�]�6x��s1%��]�[��O�MG�F��oDd?&�d�u N���PU�j���K��`�Y_�~�^zI�W�\y�qǁ9�p�c�>lݺҺ��xG���/_�����g?���<�>��3���?8o�)����[�b�U����駟�-�g_�u�s���g�����,Y�ó���IodZ%ѱ��Ww�}7�|0�s��e�$4�� ���Gq�׬Ys�=�xOSIտt��SN9�?��X�ޖ�%E�eH1S4$�p`*E'�>�9���Ъ���->�gjt����F�gX3����oQVYDHt�jL�]�.�= ��߅�=��I���BZ�cMTڱ�Y��gz�(�g-�j��(#+��"�ɓ��~���~��x�wR5jUb
S��m�Kyh<E]�K/�����'�(�����!�vt�� ���}�b�l(��F]e�R�H�~�X=�s��G���)�U�q��%Gۣy-c"�N1�,���糬�D���Q>gS!n���;!�8�,�$\�-����G�N�'������0�u��`;POK+i4J�;�����N�����K��FT^U&jlթ��<X+}�+�tzޫ�f�W��t �M�����PB) (a�u�.};''_|�E f�o�����G>�Ѓ��r����Gn��V�h�h��M�ٳ�wF�7��{�^�#i������?�|*���s�9k���h����b�k׮"�T�Kߌ��6�\�|�a���y衇.Y��SA�κu���.0���ͥ ���O�͞��,~���A9�C{J�z��V�XY��_^�h���o<��s6�ڠ:���?�c�ĆA�8l������^#�ҁ7,�n�CGqgĿ�_��O������w�������}�����H�Q#%�y���f�`C�@�C-���M�[��|x�E��h�!��o��o~y����'�C��]vf{ӦM��B �q\��J�ǥ���b�=��Q��4%3�����^�{�yzIl��O<��1o$r�����IGQ����L#:򽇑C��J�*�˗hA��J��(�K.�)|���~�����Ҩ<B�tVe��t�Ε�����?����&�N6Qw&i�>#M�"���3��尛�̓c���	!k3�x�TD��ѾqQҰ����ǭC�[�}���,����g�suU�;?{���;��E��E%�gBZN�?��>�!`���K�cZ@��~���_��W3�üy�TϨ{��_,�H�U��@[����Di�8w����}�O�c��t�;�c|5�����?޼y3�K��FkO=���n�/�̎��[��^��:/�e^��P<���G���3�+n K���K/�qd����m�A0oS�;������ի�A��iOҌ!�g�y���1����V��O%���+������٣¯j��nذ������s�=�����
�^���+>����~�R-�K�>��/��h����$=;��U=C�D�D19���Bk׮��J�d܉���?��g?�Y<��3�0�e����<j7sQܶ��6u��J�j���zzL�fi�����}�e:��c ��~E���GP�Wf=�<&�NW]'�78�y��@���e�|��LB	���X܏����Ԧ�+e:~�F�K�SLlʪ�q�,}Q=sP�T����?:g�>S��}��B+�l�:$�/�g���o�[�d������f�F�w崌�q��'��g8I�f����#\ w����-�ަ�D���.$���㿁�6ӓex�T�F��>��jo�S�@ �E��4��&ϟ?ؔ���؈�n��G.��h 8R����SN�7�)�����n�袋�z��N�I=�^u��/{𪊬{׫�c�?�����#�N}o��1���JX1HR�J�+�,�N��c�ؔ��1.�{7c��ڵ���G? ��Y�w�(�n ��?�a�F����9�Ƹg!3-"�nz*.AQ���QF�0*��_�$B/m������lŲ˯�|��y����L�xU"�U��|*�D����́,�Ȳ�3gΦܫ��Uda�O=�TF�Ӹj���6�\o��I0�YX=U8�|��7�|��� FJ���<B>��|��\� �y�>��ϡٯ|�+[�nU���EO�͊�KR�����^�=���7.��%vݟ��B:�F��d_��W����=���$@��7��W�W��-��b�Ɗ54U�s����{LBd��؆�H'��ۥ�8�Ǎ�i���4��l]m�#��=�a�lk����i3�N�j�X�F�ܹS�˃-�<z���
��j~�A���pޚ��E�ｐo���"��.����x�b�Is@*�(��Lc�	���R��g�ME�i���P�2�㱠d�y��L6�Џ��:��+�^�=S�&'�Ű�Y�f�ub����w��� F!��8B8�YH���n��:�Ro��g�R�f+�/3t�E8��G[qK�# k��+��29��0�ک�r�����`�/��!�]��:�����g\"��{���So�{�n �5�F'�l>v�S�Ì��j
��T���2�|��g�K����WaPJM�>U=4<�e0���s�y�X����x�3i�%<��E���e�����PT[�D����������_s�5����
×�8����Y���̄�d�������3�a)z���k��3����"�9�'�,���S�x,x/��n#�A�9�� �~�.�}���'!����"eD���z��i�LD�q�i��S,z��$�"x���IHEj�����$�^���{�`f�;C
-k�vO�5!�dNBo�d����"�,M�7ɢ�$̿�\YSM��ǻ���{����1��f�1վ��%�R�y(B�X�I���F�|uS2�D3+�)�=q�_V;ٺ/�p͚5y�ў�d���H��?FF�;�8a{kL�'٫�Iճ��Ã�X��q>����J	�<5�נ"w�y�W=ϛ�����ߏK��X��{U�pA]�������*Z@�č��j<x 5+~�.��!��S*���u�OJxH��rP�^e$����Z�=I�U�?�"x��K9��c���ٹc���.�ixe�O3)"���Q<���+VJ��X�j�A��HG�+B��n-e�*Cٳ$��Ё}v^�frW���*'��>z�TK桪����*�aUӍ�*��h[��E�9s��N:	4��ޗ��F��O|�g@�$�
��X��j�ꀸv�Lg�ˢ�6CMHU��d��
����1��´S�b.���o�;�a�üUh���-U�t/�W<tM�����12Յ����k���x� ���j�ׇ�j��5F�&�B������فi%�&�>ݸ�<6(�T[z�s��x��6�佌�ι�l�G\�ک���G=f�� acx�x���G a���A�ݱ�Nů���!���N�1b/�|VY�8��_�%+�h� �.Vl�V!p�-r�Bp*�+N?B_T�הG�Sp�5������A���ї^z齻vū����OZ;�\����9�k�s͹�!x?Q�T���*��3�i"�G�m��E�1�+��?��׿���{)I��#w�է��$��wD�Ud���ב�ׄ�22f�$��&�S�D��c5so%��:�Eu�Q|#e#&�e����������͜V1�>;��=��>9�9�s�=��Of��"T��E>W�cT���Z3쿚s䛎N���Ð��"=�D'��W�i��߲��������}�3�����m�7�460�� �`�$���;���S�ʘ@6�/�,U�k>�^�3�e�^�,qS�z��>�~�Z����2���ٰ��Z�I"��+�����
U������TF��g6t~��do#��u�)�xnٮ�/*c&���U5S�2�#	%��`%�L� �������=���A���HY��vѢEj��@�p�Bb��8O�̅2��w��ON)�ǫ�q�{O��,f��X�2ZF�yTZE��VeU��Y?�<F��+��v����L�M��R�iS\��-B�b4@���}8f��	\-�cq3}r�S<~����p�ಯ��5k�ǯ���w�f*A�Z�
su٥WT`T^\�^�������.\�Lij%b��,@��xG%^�7=��_t�qǾ��[E����L�6�l��'�+���h�~FUd�*[cNP��3|Ԯ�ͱ�/�)H���Ҏ�7HY@A*�r��l��!�-Թ�o����4	1s�$G�|�y�f���ձ�8�Bq	�Rk:�d#P\]�$�?%l�G��߁�nf�M�u�?)���E���� �PF�8U_� /�H�=��	<�����r��{�V�O&�z�v�s��0];��g�G��s�)�:RJ�6�O��:�b��R~��O���M7�D�)ql�>r�x
�|�S���K#�L'S����k�"�]D�G��9L���\�?��y���v��{.55=o8ଏ9�'�|���'/ϡ"5,a�ފiHuM��(6l���oΟ?��YP�m��[��\�B^�/*�?�C�2�~��ʥ�U�}�?I`�!�˼��*����$������ ��(���>�s!L��w�cl� �F � �س�s�B��2�9�8-�[*1�_�D�<J���uG�4����	����4�+��Hg�ٜӢܮ�Se�T�/�qڢ��s��!ږ�2��vU��1/�j�� {'�6��
���P� ��	��a��g� �!c�	��<�b�s�ӐGaI���N�rS��G@���f���u^u�� {\������6[�'}����}���&�]���\�*]�u����T��^�݊*E�p�{��^�
�{�~Ў��d�Nw�>�&�Ct�Q���q���v�ڵT�������y?��&�/�Q�#�#6�DUx���`ӲM��LZ��;}��	'�)LF!���$!H�C�7o���_��7�o� \(+��3]�8>��4!�e@̪U�rȢ��>Z$��c��=X% ��pZ<Ű�J͏�ժr�Ɂ�U ZKj����apU���d��jz~¡/7�L��+����U&��fEi[0��ҥK1՘�}�c��sώoq�*p/�ݒ�X��Z���b���nőZ�
�
�T^�n��04E"I8��D�y�V?(B�G�\)����xW�C��'�a	�wR�WEa$�k�Z�E�ø0���tb��'z���(:�" ��0�n�v�~P*(�`$�C<ʄ�N����L��m-C�j|8x��jl�t���$	��Y�~�2���`C.eΤ�������ƨ=�"�y��=���W]u��/�̠d�o/�[���W5�L3q��TE�5{0�M��=v���F���������>^iC��r���F�Yn�4���_]�� P�~�I'�fI���@�DW��nI6���hO3�,xs���9PrX/��"����AJ|O���zm�?Mۭe���^�x�G?���?�^�>92��i�E0/�0ݩ� 0������i�����y4��bXW�T��Zؓ����BN;U(=�[������QG�瓅0��sK_��S����X��`:���n-i������h�"T��%A�n�^��R	F,�$�UЬ�p�N˅=�9!�b��R���a���+FjU:���>[f)	u5m��~�:���}Hb�|*����c|f�J
��(���?�'h�Ӛt���\픏(����R"�ί�=Vm�I��(�J�9}b8�� �;������w�4 ����6��իW_s�5�o|�I��f^	�S�'q��)�
�R���.2#���P\�^��V�_�^:v;7:��v�AS^�Q��/uC�H.���t-y�](���-#��y�Q`��24?�p�y)���p3�U*�,��� �tȅ�i%uB~w�V���,��F{r򽧿/���w�؅v��������5˖�����m�6b��x�`1g�#�K|Rc�֩�!^ |҂f��;���c��Ο?,��M
�h� \�<��/�����&-��_�n����?���M�|�,p�RQ�V�H�jd�·`�Z��J� �V��o2ɶ�����{v���|��o��ǟ�O����7i�|r�Rj����)��V�g�����u����$�m����26$��;	i ��^f8R�т詢0��[o=�ܳ0���GjuW���N&O��ǘ��<��=i*m4y�9�����̙�1ERy��n��-]�>��@��F|i��&6Y,+]ae���mԟ$��쪷�2GKIp�pA5�1�S�6�
��r�(���X}@ ����㺯�Օ�o�+�[2Hs�sQq0���+iB>$&�}���e^��*$�_��L"��e|<5R�	���������`��h�v����� ���s���q��ݿ�vz�a�՜��O#y��$�\�����wfƏ�N�~dy.\��]�Kp��]x��s���^��tzߢ��m\W^y�޽{N>�䡡�c��ݻ�֯_��p�	���n[�f#�R�X��Je�	>�fa�F����d���;�S�������-�1.�,���W_]�lGD�x�7F'ƅx� ��.��gB��,��f��T�4uĜ*S��!@4��׾��O����x�s��}E����#���Ns�+���堳
CW��ؚ�d*>�	KD�ƨo_�V��a_Ud6����y�ҥX��k��c]J���?��칳|�_�$
���I���XՒsBxN� ��
q�pƬ�0�W0�V� � Zy(O���{s�Υ<AԶ��J.�°�vv�����jkŜ
C�ߞ�!�S$�('!,���s����������1g͋�P������ˆ٩}�L����jx�?����{��>(�100�/�7KzK��O��LK���ʢg��F���]�R�s����Zy�t�F�}4���jr�oJH�h*a�x�ӆ ʆ�ϖ=5�8��bK�8��/��bQr
T!��T.��W�ğ���O8�Ú��G̥�S!��E#:?����kxP*i5}
ӷ����/��K/mٲ��������̇��F���3θ�+�4�&%b|��ǯ_����)ވ�O|�@s�S���� ����������N˹�7�p�3��`���������Ԣ�
�S޷x���hNN���Lx�k���������`�����1�9s +��5�ܹ};묳�i��n��~�;ߖ�0^KN�
kj'�A���m�- 0=�Йg�I{��Ӂ��0�'�|�aJ�u�j҂G֛#��D��/���ݼys�^{�Ön�$˝�q�Fe$�}(i���&��u��={��f�����a�Bj
�lf�����cV��{�$��DlZ�����v(u�Ӛ�tiW��c���C����vqh��K|���{�mc�N�醠�N�\v|��t<Fb�p�5R;&�� i�`S��]썝Wu�œ�-������>�e=�ZH�WH�I�2�Wԫ��5	&PȞ�T#��i�lg�g/vF�ZN`�}�F����b@�������)7y��N:	,�O�S����⚏:�c�=��'�m(�B2聁��x/x�����~�������O?����?"Z ����̥����
	k8�Þy��*�^�$?��~VD�@�)�! �m�ݺz�j��b�8o޼m۶Ǆ�`��o|CU�;�����W���T���/N<��x��u��I+o;㽧K�X��զ���V�}�ٟ��'ு;I�:�v�Zi'3a�=a������c���:�f�߱m��rP�Z��J�4�9����Dv@3z��~����<��w�u�~;U5pkd��)�����C>~ɥ�EW7o���	��l55u�c�a&��vp�]w���o�J��1��y�%��\��ћw�}���c�3q����=�ӀG&���qS"�J'sg|��@My����?���%,�2��JC~�O�)�)�>e��B,P�������~̅S)	k��|�M7A��9sFi�ԧl.L.�EiR['?�&�w�:�J!�_"��P3�_�����=�����zi	c�K�� �d%�*��QO�k� �r��6h9*�#�C1�Zj[EbDVK&[1C�fF6
s��~Ӕ��ғO>��ll",��0h�k��h$|�,h\��5ₚ���Ԇ2[�L���^*ӕ+�3g^��l�!N�r���i�161�xn�$!8�hu0HCa�>TE�k� ���~%�t 3��/��~G DB�p'Cr�Ճ��fp���  �ݷ����JM퐅�|�=��A�r_)"i��Ï=�b�h�5��-<��S}Nz�������Y�^~�ŉ���@R���mi�)�U�{p���q�+]PGd6i�ۨ5@��=�����}e�ܶyۧ��4���ot!��^��\s��裏���?�iC-�̫�E:�`wn۱�'w�����#Z^�شI�D*�&�f�z4ޠT:,.Vi����=��7Ic����?�� �Qչ��*1�Tq/�����W^��I|Y��֭[��7+V,o6'@�{�9�&D���c�Ӌ�;�K���RI��b����d}g�*�	N�~����ıG�]��gMB�굤�9��d�Ԓ-e5�������0��b��B�hխ���f��@�Hݧŭ�D��f.�:�yFiP|����GJÕ�"Q��IC�-~�Z5��5� ~��_X���d��tCV���L�t�+�H��[.iW�c�졮��R�p��5B烼�#�S��tQq�Pg!-y1ʳZ؛S�z*��'Xfܳh�"V�R44�M�ɥV��/���������/:�с��8d�q?3~��#x�]wݵx�bb1�?�O����wܱi�&V+b�C���>�1'�j���C�����2��`xn *�gz���pq�l����*���ф9I |�7<��#/���X�y�ġ�Jm��\�ް}�v)NX�'T L�e�]�t�����}�s���.=�*ed�| ��Ik�i]ם9�1D�0�\��4��c,�������/��/_��1W�>�;�U��.�P���Sds1���ږ�`���'�;ch���8Un �U��0H��H���:��y��U?���ڻw/�b���w�C�?a�1�_̈́�d꾓�ê�?��kǬ�?���C�K��i#yMw�b�~`'��ޒ���^��ҹH��|�r�&��[㵭�!u9`U��ZXH�LdQD�ec���:*Yvײ�@gD,�����������_���_c�gP\�)Qx�;���9�s"D����Au�P�A��<�u�O��.�T��Ô\��X���Ls��F�3�l��G�g��� X���N:	��O�S�C���t����� ˏW�Z��n�	�������uC��2ď�Y�l�X�'T�"�}�������+_��9眃Q|���ƙGO���
�x������'��w |�?��È�/���0�~�V!���`\ �+���Q�Y����{�;��7�7x���;}�3�o�JLs=k$Q�{r�1���җ�t�����
(�jB5
����)2���c�����q��l05}fH��c��͜B���`�	�Nt�#�F
�3������ȿ�.&�TK��-��V�[2���(��7_~����m��F�>��]��-��-�5��K@-*��5�1r���.�%I/"/̩���g.U2��k*�z�����Q�a��:���t�V����<�������bH
�[�u���G��k�}�G4�������*����&�g�P�*J&Nr=���~�?�率ٞ>�����=}з�p�[-���C�B+
b�[[JÐR}��5���g>���x6�W�-�Ǜ�w\̶�`9�^��*M<I�﨣���@�t?�����C���|�Av�L)�֭[����v�aL+�4�\��g�cNp����J�����?l��8kғ	�ş�p�1���?�C�����o+C��{�R��]t�x���d	��� v����{�jL�<.a�c�7o&��k�RQG���?��?߽w�/�˵k�zz����\�2�̕�׉'�������l�5	�z��@#dEKI�Ase�#��fp�t�t!'b[��=�z�o~�{vS��4d�~��xH
�������ۤ
Xt�-�C<5AH%:�U��4	�0����u��y晸�g?��d=�+Y2�PS�G�'I8����~�U6��}��gV�����8u�ǰW����J�~	� �~�-nj�H��z�fnOyp����^S��7�5^c�ˉ�����[��Ά �^H]y�{���^n
��o�c������ض��e�Ӏ�)��Rퟡ���Ly��%�hz��	�>;S�/���2=Q�/% ,	�gIp^�$��HČ�Nj��Vǁo�87��%�Q��GIv��Dpf��i#��%KX��ݣz��J���?�y�ҁ��m25�l"��3� �M�4:�jd�@n�!Z���p�I��N���q@ PL��6a_����#����2�q�(ASq<�!�W�+�T��d2����� ]�.�8��F-�քg9�����(�3輂#E0�<;v� �i�>R�L�7Q��e�^֣`#~[m!L�s��7'of������⏏���;�s����PyK�!]B� ������2�+K���C4Hi�qci�>�l�/";O����^�,B��������!*Q�6���j��=At!�ka,9.V
w86Iǩ�5⻖�ė��^1DL��~�;�����������Mae����5_���{�׿��͛�Ʊ�6x��*9K�+g?&�����SV��~���l�L�����)�-�����q~O�Eq���	(�����䵓s��E~|�r�6�X�ZH�K��^��lH
A�e3Nߋ�d�蕡 {e䬚�f�؍�J�a���,EcR���UC�3u�����霘��äw�"[
�Ch�)%�F��w�ґDy��I>11%Ӥ��<*���$�y+\�8u�����:�,��rpR]�xԒ�<ۤgqM�հ��:	��m�ư{TC)�Z�l���#���g?kB���I�ߋE_�|9���EU]��#�⩧��`�Fϓ63��f�ׅ^H~�Ib!H9�+^R-�X'�x�K-  �(IDAT��?��T2����~����>��	�~)1Ad�)F�p�	h������m幡���$<brZC]�$���n��F9�mt�g����ҿ`z=�A]1':%��#��sJ<�d���-?�s�=��混n}��|W����Šeن��]�֕��
= �@�[��F�<�1*��d�����_�r~xC��N��j������<�5�ǄGQ����/.���������h�)\Uj�Fݘ���NU4�ŔRU6�)�k��z�ꛋ��z<v2hJ"=��(	 1�����!+�bqCks�̡�0��Q���#e$�706�w����@��5, ��GG-6c@��m�#Z-�f�ݒ�SCҥ������ղ�8��-�E�k 5P���A4�sv�+�JT}"A&��8��K��s� +P�[-AY�L
O���x�-�ޡ������-��:��v�h+�5HN4T�6m��`���}�RjH �{��#t���*r�e���\z饗]vg��s��I,CG�G��>�#؈ԅL����.t�T�ew��3�HN1F@�F;$�g���>�>��1�K�=�I�!� ����wgG7�&�o�A/:1Df�����(��R��G����O&a�u2�&�<iT.A{�\mw�kuT6Ӫ�#�T�0}���b�Tӭs���(;e�0�﹭�����bD�����J�*Y=ەgtQ%��8��U��c�c@�#[&�z�P�>��D�7��O�pQ�&SXP���'I��fҐ~�<��f1����k0:�+#HD	:��%!�^�� C-'�\
Ҩ���*�3F��$U�����*�Ґ����VG����U䈆*�d�J�����:����պ�Wɵ��FX��~&�R;��+�A��@���,W����x�n�
�Ů�q�>EjC"��t@���������T����Phل���@'�L�7�.u,|֗g+
2���IA�Lq� ��tKR��S*l�4JWGXv]���F��չ�=\T�f�W|g �p�t���u���+C�B%�+C.\�8���C��t�p�b%���n��}���O7`u�;�u��W���k�\X��>-e'G�����deH[с�>RI� qt����iE��2�d潊kKͪ��e%�!=�$��T&�C!m��B5,�����)3f�5���)_���z��(��/��\���.�w`¨o��3�Rk*�Ƨ���	��uQ�A[��1�Æ|�.ʤ�O�k�¶Ԛi��JC��H��&A�]?�$�x�Ŋ�y��-ߞ�#�ږ¨撗U�˲A��s���G#�2�dU
�4>�.Ԧ࿜4����NF�UA'�o�=�}�܉�����1cB0��/R�ᶉ7�m����pO�%@/���YM��i�k�B�����ٟ$TE�9����PbQ�eee����\�"q�cLJC
_y�+�EЪ�v��2$6q�e�}���ʢ���Gy#�n��3+�li�N�2���_��#X��'?�ꪫ�m�>k�,�^�ϤLb�Mu��o��OC̤�ʝ��+"$I�CO�{]?�<�b$}���$�SU���GZ��ɻ�i�f�Y�c�g�|eC�Z�(Jݚ:@��=���x,�Ow3��4dJC.f��"8�V�����Jʚ�;V2ϡR_۝,E#9Ӑ����E��Z������	�1��z��s���QD��E��B|��mG����'P;�V]�4���Ӣ|eꊐi:	�❜D��At�uPIP��B.r�eLt^��P�+�N�3�� 훊�&�u�>�"����P���Ly�t����9��~��`v��v �O�m��F��qGm�4�wC���x�{�JwxE��u1.7�x�7����;�d������1z���p��W�L�y��+T}p�Z��G�3Q�����4݄�n�~�L����ϴ�R�Qg|��$��0`��uIٓ�C��MP�z�f�@]���g�"X ��*�=��x �rl�C�rRL]L`��s�n�3\�`e��HC��2h��L�l�jHa���DL��}�k��a��E���U�bQOV�֭k�ؔ�=	q��Q@+J�4����D����i�{��R�W�D�����dI:�x�l��6H~=LL<����qD�����t_э��>���n<dޟ��n��PFX���c:�;I�m�*iuB��N|�����8p��:'�*IZ�I���Z���1V�
�+R�D�:���~m��1��R҃8��Uv���zYVjGXxe����i�H�ଯ��ʉ�	f����o@�5�SL��m���ԙ�@��u�!\�n��ޚ~sw��􌮿�M��m�\}y=6Iމ��}"���fhJ���=��5�p��^PK��n:�m���LYU��m1gZFZZݦ6?�Hӌ>��+�o�6]�1��B�I��P1�3T�~��Y�~NRj(�N�n}~�]2��U#yTK�F�C�Ѕ�.����O�vU5!ET�Fw�N�nc�p�m$/+���Ա��u��u���gQ�F$��3e#���
��d�r�:L(������w?�S�j)S���/"���,�G��fMy��M�sryB��,7u�*�;J��?���n7}X�3�����L�3f������Q����^{�={X����Z�A�����ęYJ�31��e{>��p�?w=���Ԕ�k�g0~E��sM��z�M��{8�F|�R��
	��lDQ���%�B�RUU�>$�N2�U�]U��7
���U���}H"G+z^�Z�rB��i���g2�]�{Ρ��g��ˠw!��}�ڴ����o��$���DO��Q K���e:g,H9&�HQN;8t���"U���>3�;��W�)�.�G�����iC�7a�t�w��&؟x��'���houubj�Ϫ͋����L�_�$��a��x4��!��%%��f�P>�c*�W#z��t�hNBF��{6�龦��k�xq��)k�[>Ur�A��Z_�k˖-7�t�5�\�:g�'�W!�B��2~7-����5y�]=��c�ɔ���������ϸ��B��x�{���G%V�Q�NJ��Q�E�K�HW��#��j�e�&�2�	U�rQb3�嘩Ա��9�x z,�%#�l5�P�[�zk�\PnX�-$�5P)���Y럪Ύw6��Р<���(���R�b���#Y����5�r��+S͆K�{IT0PgI�Q���gi0L��>������2�_޳]�׿�]D��`����_nh��x�4�5�A���U5*���Fz�<J,�3p~��6��{��ZHZ�Q�Z�X}�����Z���D�it��TUȓ�s^b��G����n��'^���e�\��M��.H�c����_��W_�
�9;xU[�#�Cu:Zʗ�è�4W���!���>�VR�5�O�t�A�;����L�1R��QI��h�M��E+oҀ�����e�7��E?0�Y�n�HY,��s�b���2�2eQ�H=�ܬ�����S��#Ew��2ӳP.]W���A�d��3C�	|�
�t4�6���kR!���� Z��:�JF�R)+B��/�W1�i'� �Ŧ�N`�v3�y΢B_.��&�W�����[,.�퉷S<�1a��r���9���������U�Օ����ڂΌ	�������=8=򜑼x�n�
��p������s�+X'�`M�	J�M7U�λ>f��l���K����9`��zو.�}hl)u����-�O�{�����W]uU"�
�S���c�������i�1�H�������m�����rB��������M����L�9	U2�w�U� �*�Ћ@u�����GI]A����옸�z/��v������Hҳ:R=�G�~Fq܆",���M��ο�^4�ŇAyD�Xb}�x��B�V����).�I���P_�����pZӱ8�YP����ya�8���X�:,����ԽWD�si�w�^OC�uu?H���4JШ�L��ݓ#uG���''Y����~?b�)��K|���I�>Kw"r����guD�I��04ޟO@���14h��q��?�庙*������ˆKi[;�RԱ�������ۏa�.:m$�.r��&���_��+󥳹s��+����of�F}�*FU�$��Y�A�D���tf�;R�_��z��\j6ޞ���Q�<z��U���п��+�G���]�q�O�����>��4Th��8J�5πƛ!��+B�"&-�j�������é���k\o���'��`��g�[�6F���w�u�;�u�:�|6�果l�jޟoyꩧ��\"Y��L��:����lٲ��'�<��/^l$��駟^�t顇J�'��8m?��������+��W�[ =��w�2�I�Vw�D���֖�iH�Ȗ�!�l)�wl�[�XYH�K��T�8�P�W�.aM�d�$��E^���No��Sf�r9ꙍ�*Vm��n��rb�*�񊩅�N���xCL��3�S��J{�	�By��1쀗�7���ef<P�UC>'���8p#�j#i�S+K� �ؠ;����{-�����3�����6N�G)�\��#�gR|c��l�9�%CS�V���Y����\���'��8�H΋��SS��O|f�=�|Bi'ʆ$�_W���7o���-����j���<Z�1ꩌKǮ���'>���4�,7C�����v;}Ǜ�w�\�9�m����I��AE�ˊ���V��5�Z�D«j	��1A�d�T²�*/hG�X����J��FZ��Xeؐy&֩�b��R2���<�cx'|���@�4��vlZ� �7n<�s4L��E�6�q ̅D�l߾�������d�#���/���Sj�U@�CDeC������SN9�#���0ׂ�2겔|�IOB@)��k�.��Gu�E]�
��t�9���}c�kj��aȦt�Q�	Q�����+.ohMG����O��)C9Cs�>�?ij
����d��J�&�%Q._�m�����!n\��v��],�����X�:����3ş:��\��AM��4V[q~�Ҥ$�����$HT��x�z8ݣ&ޱ���=�4�8�(��A�Nچ����U�V��L���ŀ��;:�+��l3�5U���{��|�t"_^��s��n^�����W���x���Hʦ�n �ٿ+fĆ�����m�`pK1!�^|������O�7o��~�I��??��c��w������}���&nx衇|)�3N>��+V�w��G}��d� ́C`=��ha�ڵ�g�f�%�F�W^Y������vT׽���s�+4�4�	3�؎�<�`<Őxx/)�q�Gʕ�R�ʳ�K����/����P��g��Č�l3
�A @�Hh��xNw��^��W��sE����)��>}v�a���� ��'��b�
���/��/��K/�X�d����`1DuAj�S��Ů�N�͢_�AZ���#ޱH�	H�~�z��T�����w��.�Χ"J�;w�<�s�?�|E�oGFRD�'=e�̓��1���K��/�( �"s�hp<a�)A���)��H7��W0�4+RJ�bFi�����In����§H
f7���;t��n��
��,oܶp�8e������۟��zo�e{�w��e�U���n��[?��}����[��9K�i����GI��'h� -/$�%�y+�3�l$'�f�+Uϰ�Ԝ{�^,���{0V��=�z�o�B�א�xܗ_~��_��w܁�I���RXb�zu9��8Xl89���_�,�Y>?퓖��J�7n����t&xΤ]K{?t8ֈ�·c��.͛S�q5��s��)�x�y��׿���
*�a�k	����ݻ����y晄Z@��)��zѢE��{/�/=v����ˀ������m۶��֭���6m�����]e�(`�]�����Cw�}�M7�|�� ���r����~tp��_��������w�g>����� ۳gϿ�뿢'����O�/�	�A,���;�<��񰔉|����� ��~�w�Eq�h��W_����Ǻ-��v�[��:�b�0E���Ǡ��⊳�:��/4K<�e�|u���9�brXC�W�\I�CSdupJ�${������ì�HE�R�X�kѡ4�1՟�\
��G^ޯ'�ŋ4:?�)f��z���p�^�蕔�-y��ۼ���r�>��hj�_Yy3�Y|�j�6�G_dm���g?�~��ճͦiu`�
-.��ܘ�i!H�i��|+t\�c��J�����׾v�}�����FFC�&�,3�Zl*�����T�׺�O$�Iz+2��v�?w�� �kHFM5�d�����l�N,Cr&q���Ц�M�%/?�§ӣ�M%���	�ܨ�!��M��ڊ��������~��}�������/}������x`��׮[ػw��ۿMt& }�_����7n,BYt��o�p��>������+��1�'���ۿ 0]�xq�볭�N��:�o~���! ߥW\>w���ɉ�A�����]�d�Dg
>��ρ��v�瞻֬9����/�w�=�m��n�⅛7?v��a��ǣVr׽wm~js��w�G^��i;��7*i�Ӳ��Y/9�O��޻;��>���Wq��T>�O�N�>��3@U��StV��
z~��g�Xes>0c`��K������C?��׿���5�p�B�626r����?�l�#~�#�Ι?g߾}���O�>���b���d�,��(��y�1(:_��1c��>p#�nbBn��Vp2
�XL5t��|��<� �����NpЋ/�ا��oG�LQ�\�F���A��7�De�T�.1)M��y����k<�D����=�^S|/��	�e�(y.}��p�>�]�|�W��j_�*�p�	�Ԡ	1�f���������~/̱S�ߖ�,�vn��b����W�~�?�zI�T���3�HK�$��?��?��`��1=Elb���^*q8�zW��vi#Et���ҽ�'��|���,{yv�z���`<�S���l&r%�|�*�|�͔^��D��|�������W�^}���E���@�e'_�������8����?�N �{��̦ތ�7Ə{oB,4�I�
�#����솼�v��`�}��u��Y�fA,��3N��'K�q0�Z�[�.ȧ�?���?�i�T4H\K�.*AF���LÇ���o�E��� #����]�6�iĻ�� :�bŊ�~��x��o� ϓU��c>��0%�3�<a���8��{ë� ���������.�/z�{�����3�����(��7�7�8�!pCE�ַ��������Y���J���$Z��{�z�)4��Â�Z��N��-�{�9� U��]w݅g^z�SO=?�[����?���q����H�[R%͂��c�\n2|i��}\ϾVru=qj�#�w��ê��J��OjFm�/�S��DԝNƷݫ�P�m]��wC6�Λ���Z����No��VDk������u5x���j�b�\>:��d�nNRMN&&#M�V���g��&�����bK߄Z��f����i<V��\������~�K�UuO�/g�[f6u���5"rBA�N�!��o�mh�M��+)�	��	����f��.Y��&T %`��������#G�������?H��#�= FFF��q��w|@p�y�A.�^:2rd*�B������gϙ?�;������n�ݿ������0>�B"��/���[��O2'_�p�H�-O:t �-��'̀�||��]�7���A��Y;�������wO:i�hm?~LL`<��61W��ϗL�� ۼ۝ſx���H�g[n����w�}�֭[�Ν�y��MN����-Z��ϟ?�9�g����]� /�ï���;w�lH�O=���~���Gy��V�];w����/]�v�q۶m۷�044���Hy��%������O=��B)�?��@�=��;�>�����v�5� ���`��{n+�n0L�E]�;��S�)����ɓ^UU���Hi[b�������%u۞��&xJ��}k��XɤY��Pۻ%}����E��8��HT�JHD���*SWسړ4:���z�$(eY��f��[���L�yv=��!0ĶH:�y�
�ꠋ��_��W nP�Nb�L�� _zhf���+������+�e���J;e����e۹���x��`}�?��D�$���1�[�k�O�YF�7�0�
h޴i$J_@��/�|͚5x5�+0�s�zȕ~��b��Ŵ�o����D��;v�8���da``�'?�	n��vH��v���ĝ�)��f��%�oߎ��u�ȅ��ܼy�VKX�l�G����$���6��iT���19v|˒<����0�6���` huϞ=m)������/�Ӡ���Q@g��$&ee��"�����!2�[�2�P?�裘j���c�oM����5X�_�}�� ���b��ݤ��X���N�)nbr��2/9��PL&�&?��j��ؚFOj�uQ*�X�miwSn
Y���]O�Γ�v�S���V#�T�w��\Fk{�&�=e�c�c��?�W/������w���QmT��<�#u�R/�$�}�v���+컨�'b=�CHş���"ƌ�zF/�$��%1����v˂QCk���������84�PF��U�+	��A���Q=��`���ځ���ԓr�z��X�\�M�R-M�}�<X��6X�ɩ�_4m;�Q���Ŝ��ן���<���:XI�v��o/�����w�Y�d	�k��� e�j��,���O~j�ʕ��p��n��k_��c�m~��^����'�[�uh��6�ҫ��
��(�l�����馛.�� ��7���������ڵk!�CZ��@��_�����>�F�<0�6�a�'�����|'���~��� >��&��~���o�M�}'�=�� Z����q���`��M�>��h���3�<_=��c�<��^�X���.��� �'�x��N��A#�0^���ī�'ނ�X�v˖-���/pǏ|�#�����ŀ/��H���������>�������������4�a��dtF
���%�]<3E�"&�W�T$� i.�$F�$F�K꺵�qΔe����ۊ2��*T2�'��4aYti�, ��E��qTb�Cw�)�ꏲ%���'N��F�(�d��� Wz!0�'gI=3��K��2���"ͣ'�I�/�D���1һ�CA|E[��w���Q�݀��V���ț��G۬�<�ɏ<XW�IM*�^��/\�����i��wTб��(��s"�صԈ������w��X�UƳ, w���	zx���)0Q nl�����f�9�7���t���BB|����$��h�J�N��^{��]�Nz��� h4�'�B4@��������z��n�����K/Ňs�=��^t� �Ag�i�7�?
3�6�rݺu�<� �	����W�ZEk5�� s���-]�|�_��������w0X�����S'X�z5�d�c��1
L�'>���������-�:)��ۿ��g������������#�k�M��W�����.������w13������߽�e 1~��������!8:,f�����|楗vP`�r�/�ՕrzA'�����ʜ�	8t�p�K����n֦\�H��n���:���+��)��t����J~ͭ7���5���}�����l�+�C����@e��(��Ҙ�$&0p&�T֦:��^��v8\G�9ۮ?����
��ڽ���jNc`���O�(/땵y��eD@�+B_t�e�J�W�ʺ6�>��˰y��f�*�4�,���(��/�wH�J�x��"�᧪7�-:�89���r__!�t�g�	Z���!{�縏.X�/:~�ގǼ�r�\�z?3�m����᠅ɩq����A_ejt��S׮��3��P�7���L�q�coxÕ��G���;w�����}t�q����&�˗.��O�>sH��dl u�eW�<��}���:7�p����Az�>|��=������0�c(�/[����3ItӦf߾g�����ϥ1o�޽�1��o��w��zF��������p�UW␇5_��0��\sݕW�c��$a��\sƧ�S�4_ж#.�S�,�X�
�����N[�/�?>�kL���_7o�<�����c�-|u�e�-Z�
}�/ĎR�&m��i-�MY����u�H+�?0��>��_h0�g������3s)�e> �KK,!G��Ȧ��[�X�S����xm�y�w�6ƕ���5'�a�+<��mŻ�� �#��'�%;e�k������3v���TҜ�y6�	�	W=×�[\��#S�nPFi��)A�ʆeLݝ��I�����j�-�� �O 7��}{d�օ�}̬����s�U�XB��Jq3�I&@�1���ao�+�J�5C9���	�2�R!�Ƈ�LNuZ&�?�س���A*USsnL*U~
����p��ҘY >BLs*�Y�F�)�d�@<O����31I���9@}�J�I,��oc� 4 �*C=@3���SFOg� r'x�)tb�&���|���{`;0�;����gv�Tr� .Y���F�@�Vm�,�L�.��x���}����V�� �Cg�F
�/����!������� �B�;?��9��j]�TRnț�B�n|�s�I�(��o���|W�9�ZD_�Vz�iS����Jc}�6~�{�wҞ�v��O�cA�ta�O�[����՞d�Xhb2���A�X�<�ոxѩZ�	�.Ӫ��o̅ξ�'x+��V׃��w��x�_��z���c�ꏮ�/�i��1[�����W���/�1�-�$B�<�Y[C��[ʉT�I�Ԋ���lY,;��cGg�����
��������Z�	OX�B�d�u�n��!�\
TS��L�>���g�n�\DR�ͻ����������2��8t���\��;�%�[�)9���Ƀ}�����V��뷼���2R�v &[� ����Q?�$`����anZ���2x��m���j�l�,���E	���N�;;Ϟ5-}�s��SLLy�g|��ME�o�4߾~���F�?�33�XpZ�K�bB�$Twü%1E���2YŅ0Z`�o�wo��o�}~�>F�;kxf����]��u��n�u���}T�#���{�0��J�jn�w��A�΃ѣ(s��y1���g$L΃��n^Ve�
���,�!��!%3�8�=��0ۮ���W�91��+!��.�%��2�Q9Zq�W�u.P��4���
����`B�<\R�m�2��<�
\�9����3,(�i��ݶC��(��b��Fݩ�C��E�?�n��1�����z�d:Q����m�5ڟ�u�Ҟ���ʴr�S��z��軱��3��*��4&��%�1����y\\�2���֧���H�㫕������?��O}�S)/3n��w=r)L��_�����絫�0�R$[�
��Or饗�~��D��v�m���qG�2�}�$���-�`N"$�f&��ő�"�ž}��ٽr�J���ڗ��⡇Z�x1���B��EN -W܇|�N�3�u�i�qQO��{-�*n�ԙ4�%w������Gq��i������jb[�f䕝�'��W�+��.�ȕѐZ�#�[��Z�
���^��U���m���������oş�'��}�4�r���M-_�1d�o-H���?�.k$c��R
sȧ��;5�����Wsc�ɀ∶�M����xvL+�����'��+�Ӕ��ޣ��������jG��F�i�mc����;��	�i{��JI��+��!/J��)	Ƚ��3��)�:As,ܬY�f����iF�����޽{�>]�Ҙ��?�3�4� ��؋�+�-@�l�����V4a���}6]\{���lٲٳ��$����́wP��`{i��$����=z��g�]�~='�:묳�̙�D��[(3�4��8��.n$3�CC��Fv�|;#���o���?���o��&���N������>{��*�@�~��g��D\ޤ�I���`<e�l�L5!�\�َL�ҦcLd����}�w����~��*B�9O6]���4�B�㐶Ҥ�}Y̵��s�����?'�Ξ�0v���!������v��'A{��Q��Le�w���ݤ�%��v�� ׌�,�P k*Q�̋V�'���e��мDx���%��eԜ�h���R�B���u.$/a*�i_���3a]��(��2�ז�� v/*QV�fX�d	��F̫M�KL6[��
v6��Yf��a� ;w���g�K�5��C���~�kڟ�v#e�tX����ܑ�ĳc5�ڟ�Ol9����v���u���=����T?�ȣ�R?��̝;������<����_Hڽ{7�� X����}X>�2��[n��K������>��o}o��~��׿f͚4�?�'{�B�7l�p�y���]� ��z���n�7����E]D��{x����O�:�я~�ꫯ��Mo��?>��xw�؁F�m���5�s���^"�C
�7o�J��L���pǦ����3N9唏~���:r,�*K����/?��Si������$��'�'����4?j*�@��2���-�	8'<2U�Ruq�k
ڋRo���$��xkU�%��]9*�O<�2IV%�U�vn��J�lAu���7�ݴ�9�_u%�=��:�Y�Vo���;�'*�����E���
;�{�4� ����G�󖩸zf�^/���M�g�_uֶYA������e�;�\�k��p#��LL�T��0�)pp�v&+����T���`��+��vy�豓f�z�Rl�����;�S�L��D��C�hU��QZ�d^\��v�{c+c�}��r��OceY�$���##ǰiW�Z%�N�<39 ?850��~)˵���\[ N�sgTc�R*�\��NZ�Ɲ�1�C�h�C�i�9k*�2����eں�h�/��eV�c;v�t��џ=���.��2�W������{���>8�>u��Ysg���[�8p���E�~��I���5y��������c^����V��Ȝw;O���~|�������04c��.�'��Ə�?T�)�)+7c��#��p�m��q�i'�|2&�С�����^����Oy���y�##GV��
���������޻��g������ŋ�`�����ܷ�g�^|�E2�+�xÌ�r��OI�sH�����ُF M������j�{��ۃ��<eh�P������I���ۺi�&����q��Q�0���OlF?��u���b�3�<�t�ҵk�b#��~�i��`8P�� �c�7n�10��矟����=���2 ��葧�z�<�׭[�2���~��R�`[+V��'σ}�b��"�0l���������/�r�ï��ԁ��нB�B��L���{5��ͼ�<�l�[.K}���!�@������%�HD.E�Ec���\�wT}'�[ø��k��
F$z<JҖ���L]ZEE$Q�WL����O����L�d��p�F�@I�I��BX��Z)��$�p�d�fWv'3W�3Q/g��s��*Qt}�m��O>�4D�)ۏ��-c��2�MB�&��[�T 	�+Z��u��\�5Sp������z�i���^���"��x���c��nLy�탌Uc�$�u�o�|�����R%:����o#Kw��U�W�'�9F�F�x����_�%t�؄����'�؀2��4MOj`�1�[Sz�Сm�^�`�?! bΡ�O�O�N*���p���k�Fo�,�p�?��O�򖷠�o���p�9���BKg�M��u�Y�~y��/�7��S��}�C�
 B?b�'�b�9v��Nj >�G?�0�EK=��C���w 2sޖ-[v�y���oe&�@��������k����֭[����ko�$�y�a�括��<�H�N�;��駟��ǼK(�i�-�����>���4�m۶���^�A�ٳ�}'ؼy3t�����������E����t �}��6�@6zE�?,.v���I����
�d�5��w܁�b8#�i���o�y��0W�]w����� k=+R���_�" b�(6�|�ɯ|�+����?�������ɻ�����B���������,� �+������Q(��-���Sp�;PRo\�V#���V,u!�U��}+���;]��퀆e��*�C!8�@�˗/�=}ɒe�f�������s|t��(�HPʦl��^�S����:/�ߘk�?�u��a&�i�Υ�e��>Y�b�\ P ����Зi����پ}G"����!:h���Q���:���鄪(:e�p2s'���P���!���=k�密.fWtگ^c�-�5Դޗ2
F)>�ǎJv��u�#���)O�����~���P&�xq�?��r�(�=<	���o|��-z�p�� ��R t� ��~��^4����d�Ɵ�ɟ�^�����4��f�9�,�Q*���]�r�>p`?���_A���&�u����r�10��c�[�l���ˁ�ݿ���������Ĕ�g@�����0��Y��<���I,�r����֭�ݻ伴��~�`�o�޻��|�S��N�˿����������������LQL��k ���a��	����#<�����7���O��[n������V�m�&�f/G;�����3׌3��;v��`�x��#��g(��cG����阈��@�����f�,�4�W��@�'�x��W�.4�]�v�����РtRw�S�U�Mꇊ��%�<�&Ѱ�+���"/���ؒ��_��D�t2���טs9t��<����#GG��d����w]��>�&�٭[y::�o�1�Sc�ZɲEK/�� 7W��';��/�'�b(T��R�j��j5L�eJX���o���!ؙ Jt԰s�NS�����Y}��۠�o��O��<.` �?Li�WH¶Z�`W���h�v}Dw�#�_��������Y��v���H��2�T`O�&?�m����W�����J�tH�.en w&�g�.���'���f� mA1�җ�9��߾��+?��]�8&Zƿ_�����7A�ڻw/�D!)@�瞻~�7~������G�x��+_�����6��ζ�����?�����H#/����.���@ߢf� EH��	P�Dg����|)�iRp��ƫ�	 �B��@2�}�����L�3g���C�W�X��)u4���t}�c������Xl9`1�Ûn�����߾�կB��<�x":��2 ���r�� ���30Z�ڵk��4�]�����p���/�+q�ڳ ��'�]v��[o�����Y�n7|�-�/iǿX���w�zœ��Y���g�L��w�{��W��nܸ}���׷��*�W�����%K�X.��z��EgՕ]D7�Ĝ^�J�����^S[vc�&����1yQeF�Q�ԩ�fZ��2��L�����C�|e�.0���$z��hd��E$!H<�����=��#��7�=��@0l���Z���)��GR�%���4�Cȉ1O�����y�-u��5Ч}�g������>=$
 ͊�C��C��16:N�A_)�a�͟;������h�u�[�%[X)�m滋%c�iS2ey�+f�ˤY:�,�'��-���҇Eg
�,Q�!�_�����$���1�%�-�4?��c��ǰ.ؓ7�|����������`���?�>�)H��Ï>
	�)���C̉�?�u!5S����� ��������}���� V�ܐ�f �N[�p�?8�֫����>�ն^8m���Wa�o߹�W�@H|y��ϓD<fA:|�0�zӦMP&(}�c[�n�tC��A�-�}CW1���~�X0��{��9�l\{��U!�=���>ӷ�0&���O1��ߣxoc��%�����e�9d<��������;r�嗢�W_�=4��h�ݻ��߾��GF�������;o�}�݇�m��֒K�ނuA���s |����ज़7o�4�&���9sm2h��@7���a�Ƴ)b4]V�W��t�O�Ou0��Ǥa)�WgѢE�w4�mѾx"�j�cZ	Z5]ףt*��|�+Y�}��VmOʑ_��U�8��P�R��2D�-\��D����`��ٸ��	?|iW���1̛�*�c�Ǐ=z�����T�3�5���b��C}�g�9p�&߷O���D�)��b+(��<e�
���:_[i����C#>�ћ��?���@ICm�}����~�����~��t��9���A͜&�[�2�3]i٩�X�$�w���뵟lhp���������U����	�}hkط|��E��� �`���}�z�I�4�1h���E>U��Ä�_H;^z	B�������v(�N\�p]q��~�\�bV� �����)>CF�-���z/���/�/�8�7>��� p���0t|�1��z�y�{��~@�}��;��;���Y^u��>���\�]tQ��BT|��>��ϣۘ� ��dFٖ�abD�6�zL���Rp�{��v�
L�[�փw}�� �@�@=lH�03+=���[��{���^���h�� p/�9��{hR�S���'a�u�4�uc�03��y>���T�3[�l�N�0֖-O��Xe4�g0��.x;l��|�#�����n/������!*a�� M��ح�?p�Ic@-A
�@k���~����.��^�igf�{%�$F�v���q^k�G>�r��ԟ��+ �*�(R[>��å1RW���N�[��K�=��x�7����3���/�ӟ>��LuWr����s�Ld�m�:��x��/�b^�aq�����Q7�I�Ұ��[;��졖�*뮈x"/�`i����0����W����ѝ���L�54���Cd�F�e˱�'�4[ѧ����&@7$茉��{HT-�}�?D�.c�f&�9�g]-�P�1F���qRI�W*�|N�-�!���N�T,�CUx�huS��:8iuc��$�L�\�1���T�0�x������)� ��o�+P���Ǝ������6'��>$6q��@���k��k�{�o~���10��I�B��.`σ�!6X1o|�v4ڀT�Κ�^�Xq
Dũ�+6����ŋ;zZ9��/�^����a�0R�
Bp�g�h����c�G�G�S���q��##�(��^��T�
���9�����%��{�BGw>ʤ���%�̅�A�6��!�s�=�j�7P/�z��dcD�'� �� � ���h2W��}��a�r��
�|0��~�����m�Q`��&V�A��z�{n��F��_��S�H���_ëq/ſ<U'`7��&/�ٸq#���r�-`��ȿ��^�zAS�V��i��6 9�$!s=�����Gı�he���2��>q�P�^��Z[Kz��Z�[�_Y���b�F�*b�w�+�@iF�K��/�����t&y�{ｗM�ڵkj|�F��U�{���g�Mʇ��3[��|�h����#Ǐ9Zv�}�o��	�?�
y�	���A�N��Im��'����}����Dc�,�NB�<ԃ׃vA ��>��K�t&�h�?:2�3q\��!��D�D��/�>��8,��w���T����N$S;���O�W��\[�+	��>P�N[!�чTLN1�R*>���McnBrD4��v�d��i��?���+�dbUِ)�/���������gd�ǈ��*)J��:�cF�����h��1c&�M���u�nI7�epx��Q���g�޷��G&���	D���w�x��`�68�<�P���k<8��9~�^�r%`�Cƻ@��xS@�a!����M1誫�z�;��9AO@���~�'?�IR,���{�t����rpԥy��|D�������?�3�qb&k|�Ї>�ۿ��@O��.Y����_��_G;�@��U�V0���������}<=@C~_�ւ�G��09L�K/�zC�h9`��	��i��Dcvا��h�a>y�m�C�Fg�Ba�@�"RK���E�^!վr�%�ؔ݃p���lg|<�nc��t�b�L�����aH֘���/>��s �;w�*�&��OfJ:ƾX����R,���²��I����W�x�v�K��?�i�D���Ng<�'S%�!@E>�d���������_�6<c����'��y�����_���M��ȷ+b6N�u��d7�����\$�Qj�p&y{���
�/3��qC�Y�V6 �!��j0j%�$jF�:f�@�{2и�YQ�B�0#xꀱg~�&ƼdM_㾁����2�Q��
c�i��m��:w�Z��0��xPgI�z1L\��]���u���� >R�F�13=unM�re�ή� �jZ�V�������bP�����%��|U�T�=��(੢��up�j99:Qyb�C�9���!c��b��.k ���!��S�s�����?>%H_��-�����;�.��!]iJ�	$�2Av�����>�Ŵ�@���R~*m�h @mb\5r����s���;\# 8Y)ޱZFꢋ.bo�͜y溓O=E2�$Pucs
�z��b�F��X����e#�a��w��K����Q��cM�:3<�BL¸!~���wr}C��q��6,�����_p����s[}��Λ��;A͞�ӄ�8�2m�
�MNa��x	s%��v=6��_ 	���UƧXJ�~�EK�G&r|�C;L[znۍ��ȁ�!�����I��| �u��A�p��R�X�"j����k���ހ�w0vteӦMe̩�Ή�X��^��J�zV���Ɲא�Ot�δ@�{Ǿ�~��tg?��:a�I����*�ƨ3{Lo�]%1SA��E��ߑ;���c8�>�Oq�L�鱸Ue�q����iZ�@�ܿў��(EN;EA��w�Ў�=IԐ��DD�k����4�XW^?`O�����XY�����d�Ь���;VT)�8p�q�2��X�-���X�e��&:��Z�W�3�u�&7�]���2W%��@�%�h���%��ʰc��+���N)�9�U$M�73Q���:�I�l\�Q$1��!�m�Ӕ��ô^�G��եu}��X�ɽgw4��w�����8�3�<��矿�{����VAocBG���hS�H�3'v�d��}L�����5`p���D{���e����Ҭ���+��H�n��_l(��6=��S�G�����n�`?�	�7�pF�p����!ɡ��k�ҝ�)�"H�kz)b$�}�Y��䊢L�i7Fdt�\c��[%WLsf�LK��yٽ�D�Z6����´���G����"Nj��%1I#��Y��R݉'�)����¸�
�"��&u�%g2�%�j�-���O�1#��5�c:ٷb㽤CKX>��Sf½�z�o�ּ������1�3�'�P��������`C29��י\��.U�u��_�C*�D��J�x+���Z��������@�W�B�@���[3��*WHj��E��XS�t(ǘw"EQ�B�X��?��
5F���
ʀELܚ�x75��ʉVpqFvQ$U[��vk� ���#�r��4ڰL�8��~��c�0�`�z����Ʌ��3��|���A�vI�B�|��<��/)��a��WF���/��՝f͚�!�w�O����ΧMotG�k��&d�Lq��Ux��=G8�h��
p��/��d�}r����7��:B��mذ��0/eL򗙐V����9s�PO���Ћ�"�{��l�R�[z�S��褞-ޙd�*R&V���J��@c�mf;���EӃ��o���4��W��YM�UVb�s='�gaN~(�Y��2�b���7��%����3����Z�o'�b�qj�<K�kՔ�L1�����^p�hY_�cg$�.4Y#�8��-�4�҃V�i�ʊQد�Zᩨ�oLLʑ$�~�zuc�%u�*L���r�&rz���[����L�cd�v�K�����ad�K�_.e��Bl����J#=�
�׷ȕ+��3���Љ�~*!�!v�"K�6Ń}n�5k�,Z������a�X��g�����Y�땵�Y��Ϫx��"")OL��Z��ڹ���� C��>�g~j�P��R#�YJ�f֢��+ʴ����S���=~||j|�׮=�o|����0͂^�M3��gh�d�N#x91�1(�P0A���`.h{%��xm���?H5L�޶� �>�I�A��U7- 7@�q%F��O�D��m�Ų�J7e]6W��t(فb���ݎv���ݗ�$-PS�
G�j3IG׉�p��?Ĳ]v�7H�����Sc�t�|��O5u��\��sR���c����}�'��"~iYՐ��O�k���Loέ�� 
�t�m��0U
 �Xǎ�w��<w>�t�3��mÊ�� >-N�#D�"���!�i��@mz�+Ey.��A�U>p:�lV(,$��I�XTUwb�|%�,Ƭ1�U��4��L��+=L�ᨙr19~۟�O�y��u�X^%�(u}�MsF*)E�K%�),��!�J�z�����.b4��1�/�ǥ~%-ei�+��B:�nٲE��:�3���j���g�M����4c�Ekj���<r�w��{�-]����#G���=995cp8KZ���ʠ*�S�zf2a�~*ʮ
! �� �J�����zK�.-b�O�Cy�f����M�J���ۣ+]i&e'G.����zҥ�j)qؓ1O�f�\��tұ5��-����}"跌]A�B!&��/n�4��=��\"��C�#�<����p�6H�o�
�2�D���r�3�6�ô���8�HJ�2��[�E�O��ۘ�,^A���{�ڒ��n`�7�~���t;]�=+�s����ۭ�!3��_uo��Yu�P�lI���eYV���s��M�*qӬH/���r����%$�3@����I�#wF��Ƭ�ۙn~��!D/��2Z���8('f"&��0���� \光���g�)�����=;?�\�/>��Y�y۶2��(�
�h��e1,��}��_y�fA�x�;V�X����)xp`~8��(��P��_�ˋ�t]o�����-o��Cfo�BP�L�q��1�j��Z�'�����(�����X�V����0ۣ����`�眇>1�K�)�n=OS�SS�/�X�
c�b��D�C��cu%��-%�����3:&7H�DW������]��Z6~�ϋT_���X�l����Nc=�B�-�'�Y�O�+}�o�(�j麐F�)N ���8
�la�#�8F��=�
ѩ8>�;ef�7��8��Z�7gq�uDv�9���v7گ�����Y+���Q3ǫ���y2��EQ�vƲ��IX�����,��P/VSbe�nIm��`��UU(���+&�2�?! ��RI4�$��Tk��4�L��T����	<L�6r�_!��T�2뱤RE.I7��Qa-bg�A�N��Yީ�L�eؼ���V��`��,�����zu��3Yn�Iϥ�=��N>��n�a���_��מy�Y��Y��I+�;[J�oʫ����������]����G�]�`A�c#&�W:�14`f/s�؜�Y�7��J��P�"��L���v����������M\lP�.yRҊ�8E�� :rd,���޽{�O�3{�����.X�j�*�K�Ͳ��ҊְLg��+�k�x�O�yE�9�������I%Ӕm>�4��k���]3�E�ޖm6�ޗ���R�k~�D��q�ˋn�1���2O6��EtfW�\�"6qWm9m_i�4��|ˠ$ك�jK�i�ub�I�po�D��W��^�d�K�০
�����xK�����Kb!�?��.$ˤ���!�mYقBg��ז�&n�!�E��������g��TZ?bJ���S�����jK�s��҄��_��=�3��B���N(�
g�qY�V)�teϔ�T�h ��F��\���w�q�N�K���6k��СC��k.FM}73����7����&Ǣۡ�B:� ���r��V���F-35�;\����hr��#{\NgϞ}�y�=2���w��W0T�t��C�}�v^� ݩ�< ��3��]י��:��L�;rΆs��}���4\J�x�k�&��pC�0Y)���5��r4A
��R��&�1�YR��;���^zG٩�o� ~�Cp�fE_��!���eU�$�%_J�&�11z�~H��a��YL�(\����t@�l�|E�Sv}���q�/�&(�Ȅ�CkI1�v_�V�!����2�KR��=BX���7^eW@�����^T^�6/��Das�ϩ[b�C$
��h�'L`�h�P���Y�_F�<��*QN�␕"���8Qz=V�{�х⬤��TΓC)���>������R�Y��w-���e����S$Bo�Z<0G�S]��J3+�b��X�������"z�ND�uAG�*���=LKG��	��VF�W����!-��@ɔ�X�3�<�`��@<��d�R��΀�[�}��hŴ�����S�DL���������[4�3�eunayR"'�B���V�a�4E	�L����[<��e9�r���p�^S��v���Uw)�����]���-��v?k��]���$5w1ש�Ac�MLuN�y�g.=�T|;�,B�Y��ŭ���NZ�o9r��`�%�����d0/��U�=�̶��x��+[�b1�c�V�{�i��>7���ֶ�GN$���L���Ǉ�+W�V�\�S̲ȨhXT�*�S��UA�
�fiCSTZ-�-�;YV>i�cێm���^��8Ѝ��u e�0��$�@b��9s�I�r�m&�c�x@oe*︡���r�v��5��b3�2�&ADy#�J��ì����s��2��&&��z	C^A۽��~�87�9���Wȁ��c�K���wi�)�FYV��Bi�qۏ����v��V���{�焳\�T{	��M��]�aZ0�4G8I4#$F�/l�����r��r4I�9��J�����{���$
��;I�� h�sf��1�m��y3dP�����?u�����0���x���{�(K��� C�Z�ހ�B�
��-]�t����Ś1*�F���1鋼>�מ;w.dvor9z��iE�.��,A� O����-!﷔_u�S�����,̜9�~{�)��%����ka���3yMs�Τ�}���)3��b�gQ���(�y^U m��3r	?O�ۯ��,�6��ޯ�֕�5h�z:�Ө�`�����q��w��rJz@Y���_�\��-�$��
�Sş\Ybb 5��zQ3�4����n�S�����$�pjI��Xg��ˮ�ஹ�r~��N��c%*����΋��֞ 
�\C�Q�W<"�O!��X���>^�Qzڒ�S���o�t�u�zypᣓ�gy3��ِG�TSQD?��H޴��KB�g���;�e~I���������`6��)��%i�C}��?�zdB�f�P�UIK�I"�Й��&]��bV��P���+^�e���;v6,i�/���%�ȒT�xG�N7)�+��*��ޟ�M���@+$�^��L�`�4��V�v˓r7G���㑯7/]:<s��� �{elJ���� ��	5��[�?:D��sL��1%qY*��(����T�;��W�s|5d�Z��NL0��G���_���M���xX[�Q�\�Z��֒F��ޔ���.拃��>�-��p=��y(k/U|,�i��rQ1T��n��ٙ�B{�#BT��y��>�4���VЊ�Њ\D:�3Р.�f]�9��]�q�3l�d��%�wK�H��?$A{e˪�����6��ӕ ��4���1�2��)_�%0������pZE�6b?�E����/�҉�}�E%h r�XVz����B��q��zl��q��;$(W�S��wlDB�q�>�,+Q0ڎ�&��"���Y��=�=z��7:����v ����92�,ghU��۴:�б�n�U��0���(�/X�`���t�o���@~t��I�SN�$��uF_�B�2��ϗ��Ib�]yw�3�-�I+H��"	�,�j6�N�
�����|�z�s|W7qh���F�mW�94�+.a���[�����#��i|_\|,��|�t\K5�zR;���n�w��������9s�̞�Ot]�j�f��@�J��%��Jw.5ET,h�G76��>F��/��O�����Y8k�b_g�
\��Q�b+�K�����3_1/B�LXJH��]	i6w��2
^�	Q��C�r��\_K�}�W��M�����/�jppb����sxy6�T��g023�ľS�pF)6��|:��L^ܷ�y���
'9� �nelY���J�8iJ̙�yU#���SIOe�&����w����!c�Ŗ��O��`��Хҙo)'����$=�
�]��M��fT�NݧV2��@�IH}�MxI�º�w��Sɝ�P��8�a�<z;zɭ�C{̽TQ�-��1=!���*B	ބ*�U!<����X ��v	ь9� �����
-�(��<�e [_?��gQ@`d}�/V�Ȣ�f��]���,Y����3����c���%I��&��������I.�^��>s
I�*)���@��W�����:�'?�&��4HG7�~`EG;(�Y+W�d����`�����bⵟ�$�*���:B�R�
��n��;��[L[]tZx]��/<{5k�,VN�i���D������bk*_[2�Bx�M��^os�z��ɰ�}@F+�Eo\�\�E�g~���t#�G���'+րSH��\�UKc��hO���Ť�(�t���o%�8c�r��M#��l�� Y�����Ib�i�d���h|,���0gőj��(h���4�-$�j͢&a��W4��x��T_t3W�KTEO���d^-�������hߊ���$�3�А��w��
�T��5g���S�p}��9+b>����Y$��E�1\>Dے!�췏�����@ydtdlblp�߾}۷o?��wk��)4U��S�.�e���(� Dx�駱` "��j�H��.Cc��O�A/v��?R���JT^�/y�o�Oԯ�6��Hju���yd�ES`<�*c$�_N���cD7n���5�1�4���e"T-���)�U%�Վ�9���? |ے27�"#iv��A7l?�bS�{	=����-�j���eJ�iBC�o�U�ZvQ����2�^��3�TG.\����p�~���k�sU8sK���,���Co�%[@�5�(�m]��j���-c,�Š��k6��[YK� ~_Pp�=��~T-��Ť xb������V�B���21>z��ѴQTSS�IT�9��\dRρ0	Sik��2�! �Y��Fy<�w�o+7q�e��g��md�ZR��RRoiBvR�:���$�srlu��'�\�|����� 7QЍBB�:��m	Q���!�t�hPJ*]�qd�шW�i���^�N�)8��̳���T2�J��|�s[M���-o��P{�TAK�e˖-^�زM�c���x���@�W_}��_ĝ��=�����vǪ0J�?�0S`�)�3&[(�Z�WM��SsE���v���UՉ��^V���X�jx�M+K7v��Cʬ�]�(��̫�SƝq�H��RK|���$�S�J�������5���@Zױc{02���ՙGr{�*�	jL�G]�{���"<��]FN5NP��r�͚��t�I�5Rh&͈ 2zg1�`�c�Y/k�ꚬUIє3t)3�
hF	�e71�?�V�5m�e�Yû�� F�A�5S���0�P�L��H��"��؍�D�h��4��Aq�u�����/��un�4��U^̐��Y���RNT�ߛ�"�w멆�B�S���chjϞ=[�n}��ǡ�*���?�ъM�@��0�q��� �Kr�� �2;5�YP�O��tYɦƇ-D*�\��%ţq����ܒ���l�qQszk��g�L��ޗ�47��[��ɉ���[w�YY���9vtx��v̙���%���v���E�'��� �����<H\ࡆ�K#6*���K)��R���T +���r4T��j��]fU�D�j\�K��@�1-����!$a}{?�UV��O�¢�Sx�t�9�ɥ'����+2�3$�Y� :�1v4�[!��id�	�y��t�I�8}��<f��	�N�9����g���?ݴ�2=��J+9��D����J�(A�ַ�I�l���G�U�Y��$�#��V�����F�X�P�Z�R���J/jy6*g�ɮ�h�X�ο�
���ʥ�c�9|i��J�6�� �.���ŜJ��;fB�KO�x�W��s�a��D%�2JYy���ʤ���z�S3�o�n��AeH������-��rv!c^|�ŋ-��]]���*#-�i�}�r9+����N+�/�j/��Y�w�ܹcǎ�K��1�-�	O��9c1���*�	f[�~�%ᬸ��?N022>�T�s�ǀv��V&�1)4�m��V�Z�z50�L�2��Ӯ]��ݑ���o�.��څ�tc �OVԻ��6TI�������?�<�����󑐝*�Jy�� ����_p2���,�K���%�P^�f�y�ă�� t��Q��D�i)+N`�,*~0ñ������\+}��Ә"������(���:�xV��+�ۥ�<���4-���i�����H�K��c��ut1��'�d;RKh��`�2���Zx�w�����V����33ly�����U7���#e�nnt5˪<���6v���K5H^@�X�8(��4(\�)"P4dX#����$Qw���S]7fE#+�lٲn�:%�~v&{'J�>����ʝ�	hݾ};�5	e�}�H����S]F��(3E{���֬Ys�Wl۶���S�e�g�:1���_ݳϜt������_x�ϼ%����r�=1,i�dG1�/}�Kw�y'�r<M���P��X`̖
.Ch_�ꌖ�t���;�Vԯ��x��Ě�J�W�+�4��x>��)M%�`#�n�����r����j���r:�����Ƹ�&�4l*W�%#�zY���	F`0^�K�P��5�'�Hi�ܑ'���6�%�j<#�R���ZSYx��Z2�*9Z�œ����1�Y����{��Qc���w�RO�!���d+�8$�)/��L�U�Wqę���F���PW��욶d�+̘�&�ӥ[�vI�Te/Q
�����Iܪ�4��39%
������V*��|�nA��k.r�G��� >Gx ��򘺎�	�z�7�V��G�|_��z�3/��2����m.ySK��$J���iU<7�fIlA�������%�D�ݻw�1_a�gOi:*�����H�/[�l�KپǻY�fmذ���Ʋ$Zj||�/�xʩ���x��믿��Y���Y��A��QcB��%&�"f^�����������&���OP�薶R���ג܌Tm��j`b�^hh0�j���Z4�!��O+heO�FQ�*��E�0�/�I���2����z�?�[:�O��k�;�Cm�(�ޯ��,!n�F�����W���a��ڹ��W[��j�__���دT�5-�l��|�O����}c�(tz�</>f�U��w�Ih����;{Dd����x�4��N�>\���m��X�;��k�0ͤ���?yޘI�Q���|j��U
�ݼ�w���{�SNa����&��|u��Oc=ƀDƛYY�|��'�x��� q���4p]�J�x�buq,��k�ʕ荔a����SA��<i�����ܵ{ɒ%�=��i�W_r饥ϳ<�"��(4�.������X&&sL�n���|�;ccc�
Z;q��tB����U�$�T+�X�S��2&�l@Fj��9�2�;��qZ�UQ�>-�>B�@��o^��cO/�(Ѥ��8Hj�d5�R��/rI�d�u��n�$zQ%�G������Y�	��
YJ^_�ED(�L�$'F�q�͠��v����*�qNO�\]�.��Z�
+�e�ֻ�5T+X��E�'�c�LR]�����Xd��!_j�d^3���޷�n�k�����e����i�y��A����<�ޕ�'��D�YCg�Z.�/�}����N�dm���?~IJ���RµҘ6�� S���#�܇�@�ȧ:E��<z��ϝ#��"ɺ��\B��C;	���J��#G�l޼��s�9�u�:!���P'�cI���'����rh����_�Ŏ����Wva(�n�$�:}5p��+^�3o�%�̙�q��+V�|��������j���;Fx���]�vu��n��6��5k�̞7_�E8�������B�Ѕ�ޙd���/���w�q��w��3֦��߉?oOfyB� �"�������)9���Ot��kU�2�W���<HZ+9�PJr�Ҙ\"���rc:гs�e]Z��`U`�\�VSq	�ā��,5^猄���-�"��w5,zn�8qg��>� k���g���J�Òu�s�λ�v;p�� 샽}���iFqm��,�xx��.��A`Iz��O�HR��J� �s#��Yh�km����H ��2�W-�������yPC����CT"�Ҵ.O5�R׾+�v�I;S�]<��C��X�lٲ�덜�V�7ԓĘ��x�֝�
A����v����w�y�SO=���"�V�:��w���͛7��Ot~Z��������lݺ5ϲ�����qt���6弱����(���3�\t�E�|����.ZRƔ��2YE�qddd�޽���w�L���ļ�t�1]C*.�I��Z�V9?�������Q�z���
�P״�Ӌ����uv������/aV�]X�	�"N��as|����yҗ2����H�^���Y�RNS�">�+i������5��Ͻ"3Q:'�۬1�A����3L�4 y3w;S�F���Y��,�Q�|)$sd��hS�&<�Y��I��33S�D:�-�D��n���%HB�sgڎ����f���M�a���c�o��T�O�hS��i9�S�-�W�`�c�2dG1��a���qQ�FlϫɌzv�b��/O� M���Re���O��^��f?�fI��cB�[B@c
̼�%��<�û��1p�u�-[�H:�#c�� :4~Ю*e�>�e���o�뮻��y��z�o�A�,�G_樚9sx��gϞ�T)�\�CӐ�!b���EC��81Y���=��_y�������G�~r�g���kׯ_�t*�w��a?����{�S?���c�h���ϊ�j����#G��T��zv'���Ai��҅�E�H�H��!z-Խdg�z��-q�q+���~�LZ�V��[$�q����V�B���AZ�h��u��X;�V~��Pg2IaP��}��1�P�;uk0�6���
��a����u^X̀>��+KB��^+���t!�q���L�$�^`e;�{�th*%%$�jx-J?�@��
��b�$24s�l�PC(ya~y�%ָ�v�W
���E��rzw);�p��<L��V:�c6����ڥ�TM�s��s����z.*�������#GV��A�1i׆�]�N����w�I�_��Itb�(0�ﭷފW��W�y�C3˘zG�L�:ؾ�RS���ʉ���{������瞃���3f�p�v�^]|�Ő}�̝NxϜ9s �+W���Z̷	��C�ݫ�����&z0c�0F;15L�>}�O195ՒPu_�7I~��'��9�ѝq�C�������m^p*';tG+O햾�5S��!��������|p�O#����2�"�J��d1Ȫ�TṰ�SƳ]5m+Y��E�6E.¨�n�c���$������Q�+C,�ϒ��G����H�b@M�n@�� �I��{�)��O�%FpPM�#pP�rJj��n�_���T�(厨We��!J�������q/)xk2�`|Zc8�aٹ�(p*���1�a����!J�F[�����|�� �j�Ǫ�������FYT�����Z�� [���%֧��|0�%�[���0<��@�S�p�*S��ʤI��J��N`��vz�ߴ�K��<��(�^�n��!*�[�dCj+�*���9�s_T�����$V$����Q��W\�q{*M[�̖�0��rM
bT�� $sg�!fb�O��d���C#Ǐ��<�O�e>ՙ�$p�)�a�Uu���cP�O�3�6�����[�;ch���}����n{��K/����_�f�@�K�|����P���{�P�}3��8�ǓO<���}�=�}���+ewhp(KZg�u��� K���Jn�SNY�d�[��1�*��1�ŋ��-o��|����R���� �/N+��� u|ԧbٵk1+Ӻ�>�L��:���q6 �Yص:r�h&��4 �TG����>_�F�y��X@��EC[�Q��	��py̕�b�)�&����*H�|���SQ�4��]t�*����s��-᪅NYK[R�籴f���eCCd���^��#b�^���4q�������-�*R��G��v�D��E����pTK7�B���A.�S'uaM�)%�!�15�,:Si��ї��;��@�X2P�H�&���6�������_��C��:��_��U��ߎ�l��Ox��Wk�Ό�m�^i��FN-߮���A�C+��n"��i�B�u�#�0Z#I~�2�� 5���ٳ�CF�gUxp�������4�0Rĉg�֭[�o���O^r�%6��j�*�p$��J
��n߾}x����z�����KE������d.<��k���g�?��s�?hu�y,�9�1i~�Z��e˖]w�uh��?�1A���3\H����d ���>is)�z.�&��E����dɮ0N 2}IY��DA��v�T>,���>t�PKP�)�+�?�5��ќ��2��/��(;Ӎ��'�aM��1B!�0���-Ǝc�@j�����!��4`(+�r����;�=�.�Ӊ�ajn=?����*(qQ�e��m�Ob/�أ)��_{,T1�1	bn�'Z�I�5Fg8�6�$Vڶf��;��G����	�F��i�Q���;�k�WW-��^�S��2cG�PjV�9�NL���S�zd����E|K��F�zZ���C-oV~jL�o�.�4�f�p�E����ehk�۲�U!���Da��-�K�w61����S��0���*#,Ġ��0�V&��j��� ��G��|C����:t�p_���e���~����L�}\��bgjs��V��ݼs)�[PX�V�WH�#�������t�On8g��u�6l� ~�� x�t�?~|��͏?��� �-:'�:�29:u���W_}5�|��w:|`h�o��y��,Y�h��ӒR�6�����N�pO���'���̙â��$jIV�D��ܥ�<�[��Jc.J�J�*:�r�[����7o�ƍ1�:.��d����"W�ڱc�^yȐ��d4A�c���R�N�M��4���,F������y�mFI�N�����Ջ����Ϲs�ȅ�H]8��c:����"��McQ;O?T/q�wMwic�cLPqտ")�Q�w�)����䩾)?d*d�FL�¨�~
�e���)��؋����21�uj�W��Y�Z+S��U��6��%�W^�}U�ۤf�h�C��'�G��8�_��t�����x�`o�u�"���g�ISw���ۙ�Ҟ�������0�B�?a� -�Z��֔xQ��n��T�����ŀ{�JN,�]ɑ�ϐL�ϟO��~LL�W"W:g�����2�4Z�J��}!K��lڴi�ʕЧ��c4����7���m����N�:o_|�7�0:v�s������*x�>tꩧ�X�B]M�jY)F��իW�|������{�1 7e��w9�lʅɚO�m�Y��ȓ��bM�2FrO�aw"Y>|F$i*��Yx�C�d���]�\StE�����M%���%dǲX��xԕ�S��9)�E�'D��	�[~�}�ȧ1%u��8�r�H���4��21������S7�>/c�-�G�okb\���l��'�~\�s'��R��2<L1'��̤���ޓ���tl�/�7;.�dY��E�R�){_w�E�,S�J�(} ���\U�[ƛҊZ����-��9^M�U[��O��W�����v�\�r�i���Z�`$'6e�ͺq�yn��v�>_��sW1�L�]ͲOd��[�\�1��8�<��S\�b�c�6;�$�&T����nw
S�jts76V�7�-���yby����ޙ��u]w�U��{`7��(R�e���H6`(�^�"��
�J^y�l���$v 3�I�Y!��Hʜű�lv�������߻�nUӲ׉�����p�����ՁX��w'&��˗�\�z��y�(4�kc#� QkApnf��7�|��w�c��/������+�{ݹs������v.,��T�U�n�F�q&#߷o_eٔj;���9ϭ�%X��O.�{2����z����G���]��6P�5tme�=�d�T��3K��կN�|�?�����O��"X<i��֍�A�x悇�����bE�빹9V��t���q)NLN|� b�ېh�&�醓&-�d�[ճh%w���]$�9)�X$G(�x�*��S�z�q�P����q��2�N���W��p4�+cz_ZFRpBO � ֝p4)G�>6��\�J�ɴ�a��R>b�o����������"�Y 8U��{�s�w>�j ��H��W'5 �X6:���4�}��v��ސ>���אָܱv�����3��Vl�vr�wu�I�6gertk;��
n� C9~,�@x֓�A���L���\�ԑRG��F�	�u'-��m����Em��!ޕU�1����
�u�����3g�H0�L�b�`���_���Ǐ;v����c+�b��,��N��e�|������\ȧ�eդ���t���y�1�fft��p?3�Z�"4%͂�n� ���
ɶ^���������S�N�f��#~ ��8�鄡�,}��ݾ}j��H��sp#jʤ��A��.]ڳg������h�p�g����:7X�^V��.[j�i$&T�VĢ�`�֝zQfl�����¯8iQ��&_�]mfV�@�Y-3�F���QU7Z��md�],1X���Sj\���w���0J� �y���T�T����ӋQ�I�|�6� �`}�=�Ʃ���سf�kr�4M��Af˗��|�=Lh��̘�5�N�@0�Etᤨ�%v�1HM�L��ץc����2c��T+n��(S�����y�� �+�GT�<��6�mz3^�+K�`��u����
4�%�*s3f16I�/��JP�'&�EmD��);��㺦}O��|c}S4ӝ��Χy]���o�9�L��D�.3��K�����+x/�Z�������z1�c�;Y��O�ٳ4?��n���ɥ]�u� 7�^��8�cR4�'NP�K����߸q�]�E�w��[��p�������i3�c(f���4_�i���a��9`�e�t�`�'?�	h��x�(�X ����ͻ���j��=z�hee��?�����ڵ�޽{e�`N,Qs��g�i��P=�`ka� >p�2�?p�����K8{��]5�/�ܹ��Ni#-�����uuu�\�Fz��^@��ݺuKKP[5iz�W_}%�O6	h�Z=$�G�@���?�TbTt�F�.i5�~���������L�h�׺��ں�g-[&Q7��Q�{0�ܒ�_��~j��3!��EP������m�,�o�:���c=_ǻV,?��=��֠����7�[���b�m�[(���yn{l�5��ӸW�1�s)���]�h\r)g�x�j�X��8�'�i6j��7Z�A�O����~,1Z��0��z��p]N��z�)�29����m�)��Lk��a�v��p�/���>Ì�$$j����UT}����^{��W�U=l�J��c�S�Ol�ؚZ6��ɫl��67��L�ZC��k�X�R���K;T��ڀ����>��b�����3ڳG��w�s���*D��$�e˩ħ�Zo�@����(����ϯ}y�Ր~h���!������Fi[���jC�u �d�@�i;���͵���b�[}!|��~�MI�.|�_�����ACj�I�ۖ��P�
y�2��;w����~�i�����q`��׮]M�np�re9�Ԏ���|�8���ƺ�G�������P� t�7Q4ز�!,����4İ��z��3.��H|�K�ܚ]ZrF�Wc���;v�e1��U}�w׮E��OM�2�3�/�$#���(>ԃ�م�^Od'.�F�� ���"#�ޢ��vJXģ����z�g���j���1m6V<�0MVA��=����b�
�~]�����E�4z)*WG�w�EL������f�g՚VM��Z3�o���~��}z;�Qh��g⩬�'�М��`Eo&vH?i����jS�U#�7\!*���h�{5�X�@O;p�����=�c�7�_�9�#n�o���2���<M�v�̚�AC'p��q�TvG;H��9���~
���%��x�A���	�͆�2� fL%s�����+��~��ؿ�e'���v.,H/�D�����6A܁'��97?�A��a{s�e�Q����zC�'T����CѼ��zf�����/^�^^{�Ho�1�Q#�nga�N{f��#o����}Yݶ��p��¹��Lħ� ��������F"̶��.ASX��Y�o��X�ޠ����W�����l�1��������~v��%M5�X*����b�S9�g:�q����]� mE}#j8v�ؕ+W(�QD�����k���+�ԉ���ꜟ yX9��gB� 1���<�)��G���{?��R0��`�t�S��"�곚����7�߄0�n��L:d��=�偷�[��>��{Ğ1q������6|���~U0cbi�e�X��R}��d71���ϟ���Xk�vߎe�;�2�_����m�F�BWt�HW��WWW���4-�hQ4J7��0*`]eT*ٴCH̓���2���Lύ%l�k���S��y������K+�u�X#��v���q��-^��ը��X
�̚�t�E`���4t�5ry�V������M��$�r����۲���/�����E�,4"K��LO
��14���efZ���T��o�Ѷi|뭷����-K����ѣ� V@0pw'��D0jJ(�ݔYr�4�8#Ymnf�>0?���-��dcυ�Uq�.����*��%a,,vm�]=(�Yq�0�2�h�8�I����K¬&H��h��kWn޼�I����8�ik4� 7u����ލ�Tc�|h����~ }�AA�L ���A.n%��+h�Y����JRGA�84Z�#�i�ĵ���'H�⤗/_FJ����zf:Qs�¬T����,l q�H�pe��U�~T�I5M�-����$�aT�X4]���f)�qߎ�� z_K�QWP���s?;�*�٠����^-���2RBS���O${d����4tD���Zϝ��*e�鐕0�i5Y_Gp���q.��SQ����={��|>����lm2�&殔ܺ{;�k33anm\�2K?��,��;7|�!���TUè�S����[D��� �	�	���u��rK� b�����'�g��$����N;uv�܅��~�׍K��QCj��1��Y<�6�t��~�"Nus�X�ci+��9�w:�b���� Ҩ~���?�!fC|E4��7�8-�k �|��Z����������G+k�֯~q]K�|m����{���
m�y�b�ذڑ���rA��w��7�����YUoI�������PAC����FD ����;wn�JM�����Z\���!d���G�v���;y�ĩ,<|�$�ux��`d()}`=��'Q��ի�ҰsV�r*$�S���Q&�4�@暘��7���mj�@����C�l"�h����и�c�1��n@��Ckl6OȖ�9��yi�5@���>D0�A���]uS%1��(����|]s(�#C!
f�ҫk�=����R"xO@7'��g�\�Z��P�1+sT�(�Ρ��o��(�q$eP�9��^G�^#au�
��b�{A�����K�hk2&BܔuW�(�H�j�,�.p�BlU�h��[��{��dݳ|i�Sdv���7�F��1lIMt��9п����I�łƠv?�Y��bVMԳ)8�d ���AW�{b���P&���3P��F��0�����J%���[��#����GM��:E�:��c��c�A �U�Լ^�R��Ϟ=�c ؊��tNS]�r�W(�������B-� ���g�$����K���4*���)I�pPxgX)��0޼���ɓ����$ۈJ3D�s���� �]�5c(8�������_=qJ�1�h"j^��'������33Ą��K������7ߒ���_^��yָ�[+��ܹs'D&t&&�����D���	U�$<�OGO�A�J�T��BJg�j2u��<�U��7l��$²r0:�54#������A�=�!�9��ӹ �f�x��2:�9�cfj&$y�,�=@��Q����rJ3� <
���3�D�+f�	vd�����e�� ��9���q2R��*�3�S;��n�e�'3��*yZ�(5��?rGC��^���~�f֢c\iʼ��m�`<]{��2u!�hY�<�֥���S�g&���	��g[�f�c�[D]\��ۨ�,�cV;�2�n�ϡ:@�z�8���ǩ�KL#:��=\!�?Qn )>��*X\��� hGR���LSI9K\��X��!���|Q%񣩹2Ej��V�r���=�q3M���dl���P��h�f�����O�j��"�Pbi� \�:�CX�2,�
s�b9<������ǖŀgb��l��V�纲
�,܃���ǐs��U������;�2I(�qB3����J�س�p��2D�R4�s�J]�@��jp��g����*d�+BU��W6�ez�U=��V���	�w.���C4� p�N�޼yk=���Qpk���y��rz,��k��,
�u<��7�@wc�[*���#ݴ��A�������&�:C��l�D�E��0����� �Knf&ٱ-ݸ�nH~	��;��y��������M�q�H��N��(���W>�B́9 ?��3��n�}��D��U,%��{��"Z2|����F��4�\.�G��A�#DB,ͱcǖ���3�;ٽ�(�A~��Y����|��Am���s�fu��_|�l�����a:Իp�k>�t��ùo��*L�X�kN,F��a�YԦ�+��[(Ŋ��3W�A��Q����T����s؞[{q6H��hu�$`��R��F����R��2&SC�w�ߎ�hrJ����^�;]A/��V'�9�z��a�yGa�!v�;�g�mD�����׺��`� ����K;�B� �<<�/��4�l�M��phT6)�m�C�>\D$q��Q]�y���	oː���:Ir�2�mf�m��m1���PD-��X@cO�"l�N��E��׎>ur��F��UƊ��z���P�jl��@c�U�G��R����4U��b�/|�ԓEɫ���-;N��@=�%�	t3H
s���8����BA3���xT��Ӟ^
쨢-zx�����������χĥP�����=|�P����;Q���^�Q9]j�@_H}��%�j��'Ooܸ��LM	f3�buu�ƍ[pa�ѣ��ٳ���@�@$��p�s܅p�!sf�9���n�\�������/CN�-��Z?u���	���q���O[����(��f�^#��!��I�����u9Ϊ)RŨ���a�޽��-`����a�P
�߿��O�:��M�_?~,NC�#��G��򜝘-�Jv�ǝ�:�̃L<���L�e����K���d1Zm��me?	�n�sv~a�uh.Z띘��9T�v��]�դ�
�@��żcU�!�D���ʜ�K��:��dǥOW�ø�c�Y��Ǹ$�"(m�Y�����/�Vߢ�9*�ڙ�.k�Q��ؿ������=�G�/��}tiiif�|Hb��!�R�Y2���/��Y�"	{t��I�7Lհ�bxB��t^m���ى k|d�"�?��}�*�2�������~�ّ�O7��[�W�j=zY�:O���F�k�-�4}��1\:n�#�i;��zPQ�2� ��$b�ZQ�T�����?�?���C��������O��W�^\^�pA{��������{��E|�B�v�x�L�h���_y��,XA��� 8?��Z>q��ɓ'������k�3lB̩j����ǿ�����Ν;����,I�m��p
�����d�����0Q��8vT�S�0z�&�P����o>|��!~�W�ݻwi�B@t,�ȹ�E���im(������]k5�G7tϡC�$n��꫅e��{=�F��«پx��W�F�9sF�kf.]�$N	�����V�>�{u��A��͛�&g�)�Ty6� 7��s*���uj�� �8l�vr��y��a��rՖ1@E�1��]�a�8c]uN]�Ռ��9���D$�Owz;v���D��,�S�b�:�(o5f"������r͉	i��x�~=���l����^�l��G׹�Z�,F���vP�%�,���?��@���lr
N� ��Yk<�|���YS/ˆ.�54k�g�6���byo�,������
�f�<$~m>47y-�m���ö�7��c⎯���o��g_Q���i�d����i��4���8��U����Y��@����Dwjjz����U�����\�n1In�u��3$��2Tiԑ"�q�7�_ف���@�t��A-s���Z޷�����L�D}?�K�<x��գ���79����w.��1c���{���NNWu~���F8jw�"�1)����._�����|Er��p%���{����a�l�XJc�Z%djP�,ֵ��?��������)bn�{����g��d=�Zơ
;w?'V,.L4!�z�s�؉3�]&�YnK>�v9��G/W���4r��`��R���QWCYk"����*I(VGK�k�髳D0C�^�v,,!J��,�)�m'�x��^6�K*���d8�/6�(�6�B���'������ٸ�4ݛ�)���K!�E�U���Nu��?`h�6<(4�����N�g����¡�����Ž0�,h�۬	�b�˰�O��_��W�ad���"������N����r�c��-�E��1���z�1�a��U�YIj'�H�q�,��n��A�DM +��fI�W7sI`ĳ��ͭ$��Oc�! ��K��������D�A��՚P����<��7ȝp_ef�	K�bo��=�4�O�Z?	�%�zdgC#R51��T2�˘�*��N�ĳ�yTU1�`>ʌ�8=�W�nq�PE�_�M�j6�Y��<*���}ғ��[�s	�B�����@:p�wcl�$\3)BV4�����D��v��靟��.;y�U��Vͬ�s���Y����y6��|��W��q���<��Ε�y�/�DI�35m�E�Y�N�.w�N�c��:�ϙ�t6J�uL�z���0U¹Dy����eIඹgj�-��G���`��K��d��� �:C��"9m�3�֤vLm��0��X�wn�5����S�0]��c�V'Be+���f�T�N�x��H�pl��DV(^Vx7}�?�f��>^���|��u�¥;�!%]�s�����0����&)�+˧��%���0gf���dPY�Xݮb��|���g��X�qu��Lc    IEND�B`�PK
     �;\ŏjY�-  �-  /   images/f78ae6cb-3b21-49f8-a0a0-4b83f9561715.png�PNG

   IHDR   d   ?   ���7   	pHYs  �  ��+  -GIDATx�]|�\�uޫ���l/��.:@�$�Q"@le��|�gG��H�?�b���gӉh;�d)�MSq>S�M�$�& �� �(`{/��g^��}�v�!���y�{�=�?�)w5�u%Ir��?���c�,��{Y�]~�i�{��F��vnn����.ˊ��JYQdIrUU��e)�"I2��]|�(��^��~u�SUŶ��.\+&�_���M�Ę��v*����l��l���з�}ըX������F/]�18�A��rSS�'N�%��4�mW�8�P��C�����6^���O<��C2hz�X,W�X�s���|�T�.P7l�+��i9.��h�.]*I���|\z�$>�,ۖ���r�F�$�?���-����.n��\�._��H����Q\��既8t-]���
�$�~��jQ}��w�F1$��ܔ�ƣ���0�x��7�}��o|��p�ֳ�>��3Ϭ��E�F���ٶ�-��,��#Ɋa�@ 	��uH�u�T*�1�d��gK�BK�j�dQ����$�i�cROJ�,,J�&�Ss����X����{�u�d�6���?��Q���N�:|���t_�JCͱ@��[�NGCj,4��lٲ#?��s����=�	�Z�>��O�ᐦH���C���C�l6���7�|����R�=�b\
aAR/�����<o�Ӷݺ�ԁZ[[yI�\p��F�vb����V3�5�]����-̭�<ۄh��%��� DP�t�w۩\`�Rs��2�H@����D�OEnjj�������w�{��?�ǲa��g?�������fgg�'��1����w~�?Ij�T�ԥ�{{{�]�Ǥ04���`�u����MNN�HG�KU�x,鸶���
^0M���Үj����-��QX
������E���鸬�nMOa�|Y�Kҁh$�v�QH^ޣ��� 	}�J��.]`�S�O=�ݝ݆	����p8~���<��9�	�\.cr�*��{ko�\��6�` �?kH�o;m>f�6�7�{���/��, �	�BHP��a�0�x<N�`��Wss^�rey9���Ė%���g����F�0V��C�<�ɉ���d(b�.۴�^��&��wi~,�e�d5�����M���.&l544tw��`K�Z����'�[��`Ld�FՐ\�Ď���S�{�72:*v��䚗��at��w��ȑ;6�:uC���b�d+�~��h�#�1��~��t:�9�>}zaa�7~�jT124tu�4�;�h5M�M�݂�C��o�طoߚ5kw������×��8����ۦ�s�!� �$�J�W���b�R�5}td<����c���X,v����̢� Vt=?��繟�жf�M7�m�����o��&{.�J� ��ѱ�
˻p�b��7�]3MK萴�X���e�-���2�(� �A�4U����,��C@�R��8��_��J�:�t�������n�]���ٽg7���U���udb� �� p%��z؇i���}w�P�2C�0������������͛�@��?��Oɀ���{�B����㏿����LNM�;@��)'��[��?������W��Dc����O�/��
:��H��y�ݭ[������J,�o��z�7<<b����C������ҥ� =���&
q���	H���=�7
; |U�VeAhd6>t��	��C��Y�`KI� ����j$�-���"�_����:@=�/ʒ���2ۤ���Y�,T�r�T~��n��d2�I]^�׻~��J��/,ˊ��U&��i�+�6a��HD���tSc+�P(T*��
�	Z�&ܮ o�bB篾&�OJ���dT���n(��GGG�O'�l�^m���~�W^I$�B���Qdj/Ӳ�S4>��๩�Y 
�$��e��M�6|���a�҆� xp����k�v�K��{���\�����2�����R,����>�y���ض��h�j����@��V�n�>w�Zy�Y /�����Y�'��l'.q=�L�_����ԇ~�%�8ǣ}�,LZp_�*�
�
QD�T4M#&�	!G�L����$l���J��a�<�AQ�O	�!%¬�dR�t�t Dׯ������pl�EH644�n]�X��L����$�@�1-A��O�!H���M�d$��x�=
�Úk
o����G}�;��Ι�g�[4�����F�Vf���ߍ�H��0[�R)���Jki)��Ӌ'NOOC@�����R6M�^�&-���%��!H?��D,r9z��Ç�z�7fsˈ"0r.��w��:p����x�~>B}����g����J2�0_��0P^��Fm��/}����sg�0�~U ��h�	��!�E
,@M@�Tm�ƍdkl.�im�#�p�w�ҥ�;w����c��oim<~���D��|���?02r#�+�����۷��E�a(B�d]ld�Z[{۩�e��bp���ׇ�����8�7�ܹ��ݻ�P`�
U�wG��v$�gc�X-`�ȫ�b��ea�@`�~��/~�w���W'�BJ��P/�n��޽ƪV\+"�/-�H��� DpL�BX.��M�B���l۾=��������J���C��]*��[�nO��snٲ��Tl�loo����K�>�����O~�S��C��OkR��Gq�@�������AH�W+���zf	��H�Ӫ�A�iy4��@@}��:�_��f��ڕ�t����*������؈1m��Y�}��P�E3q($�6_�~=U���/]��s箱�( qii�RKsˆO�9iYL	S[\\e	���U���ڡ5p���F��x"z��U�%ٞ���fs�m�"A[{z��ZΣ��$���	��̖��S��#;A�������K�R��ޙ��]Z��d!STg�;`1"&3&�U"ш�r���33K�yB�Ca�#A��&`~`�z`ΦX,���F�/\�D�}} i���;�\����S>���:8�$��5R�>��U�!���7SASn�i����<6��!�x/�-�l�C���#�Wy��Q��ae��2��D�59��_V�I�섪��_6J�2l{I،e�? v��jsSS>�C�-J���LwC����{o��˃�m�D�g��t����+�QU�d\2p
3@��0qD?�Bpi=@�5�X ,Xv)��9�~�n����q��"����AW.�D�e�>*�kg߱����-�CFU��RHwԀ�Y�gE��H[��)+�� �Ԗs�IZPqE�>rmqaq˖�0�b� #�J�,��}E�|�Ro�Z��3gN�H!�` x�����ɛoށ�jbb���R^X^��o�J._��'0B<d--����_;`$*ζ�딇��8uQ�M�65R��#��&"Q��a�O�O	��h�����*e`rv
�z	QDKg��͙?P*�l�"��~�ߤ��wO����t������@�t}z9�mnn�������e2��:	����j����p��y˶��^�嶃�����ܙ���f��q�� E ~���Ru�����EBI�$�J��1r۔Mc��DZ�Ҷ��I�@��J��e�H��V��G��HبXҲ�,9�%e�&5���<��
��=�d*mA	!��I$b �жb�"�ה{�{�Ě5r4�O6���Ҏ�;�f9�L@�;�k�өz�oX_��Kѻ �崏57;JELB����P�U�#RI��ֵ�	�1��x䀳*�GW�j����{�Z�bm+�*��-[AU
 Fv4��C��pH�Tʔ�:�Ǳ�1 3��v��-�Yf�ncC#��\-��ɺ$�x2Qw��w�m*18���S�����%+F	OX\X�4=�ҍ0.A�^!~��G��UD�����oD�z�`v9���2X�c�H�3OWr�̵��Wb�J�R>WP8�Y�J�Xd
ULմ̏�(W�&��f���|U��Fc���s]�s޲�ڶ��+`ʐY���!x���Hdx��XWgwg������lyqa��c��[���5]���#��R�՘"��u�SS�>��\.��]jik 0�uC �jŬ��]d�(����a��y�V[]�`b׮]۷n�{��c�|q�����{��K���EHP�V��͠l�d��ϴK�Sue�j��	̉v�ٮ�U�����A���U+���R��N$� ���3���m�R1�����L�)�wR���ա�]�kLӶ�v<G�I��(=0t�ں���77����'��2��Ƙ���c�_��j���B1���۷Vk���)Ѫr�j�E���
Kܶu�7�DSS#����C�p�����erz��kf!rɖ���ӳ�I�aM	�ZS�?�V,_���<�tD]J�r���L��Z��ӷֱ(7ID(%�H��߇KeWh(�캺���8��t�ÎIӡ,՛w� ߸������^M@4�v���Jn�5�2Ŝb3�Z*ɮ�IyU&F0�0^��HǏ��ݟX\Z��j���W��Vel|�&��2W�
c�r�t,UV-�U��Y���R���-RV%3V+�,�9���9C�,K�w$�/�A��Q��ت)�E�P��J �� �St�"6ю ��%KB�ɐ�"Q���➭�A�%�Me$��q)��z��
�4���W�|Eԃ�kW�=�����2`a�H�� |�T6�fU�hq��t<�⤷��Ym�BR^-��5�خ�!e2��]��:�"����N3K&��A	m. W��s�cs$�����
���%��Н��j"����yh�\���O�Bp+d�khG�T����Q  NS-'&�8�s>�Y��Cz��t�-EL�/�Q���p³}��Rr��\�����Q~�inq�j��t����ή[�&4:1Tƕ�#�@}�+��c�m�4g�f!�t�����-��X���LSs3������u]X\��B�B"�'c���F]&�4��J�!���"3���2�;3tꓲڜ!�����7����}���陹��|��.�?��˯\��*3TY/h;�:!,��+�L	�Z����v q�F�D	��R�,~�����dwW�����x,��-�x����"ȪY����^�~mÆ�
p�p�����d2mm���ZZ[[��/�ڵ;?x��o]B�_�x�nH#V���nlj��<w��m�o�h��[�m�p�!�*yf(�)���wll��N7��O#��b�;:�Z�]'�vW�!�[�r�Z�n���4= �Wj�D�g��lb��5�\ES��g#�`C�!_�#��hm3��]X�a�ajrj���� ��݃`hvn,��T.c|0����l� 6||�;&��|)��Pj�����!Ǚ����~�6ggf7�߀�tia���)���ժ�5��������z����E({ <��_��ؤK�/k�N��� O�t����6��	hN$��R��8�V�x�Cp>�@M�G(��9ȅ�y�0�8;?�G�*5��C��_�űI��2g#��ɉ��V�<51�F��K�~E�\�aq��0o�ڎ�n��F�G�[���@�q=H�<BEӎG�UӘ[���섪��`WVM����Z2�4kzz�{�� R׵陙�ү6�88rW�Ҋi-պ��E#@b�ES�L�IVV�;�U�������ծ�f� �l�����`.۷[�;:6�~�_���ѱ5�k �7F'�d$�./kjR.����͛�@.�����&�^���V	������Ucq~a��uϰJ�l@����E�Q��8]�~�먡�i|Ϯ��l����m!V�i�6�����9�е*�Εʔ�sE�v$%�qG���N��{���_��	֨Ϡ���l6��"���(��e=��ض<�O7�Z�[�ojf
6�;���q�@hiy#���J��X�n�c��뇔/�#D��s�3�2���R&�q�F�6�ǆ��܃������{#��o��]���������^��1ɫCW�k�C< 2Q��O�� ��*�%��-eM�sj�-�SǒSK_�G��Z�����3r�w���6(BSs�h<�i�F۱\�AlA!��n޺�]��~`=��i677� ��޴i��:]w�ͻt���u}:�ĵ��TsK�?B�]�w	z��U]�$��D�ʅ�uG�?Q��фz�4��R(H$��Qikm�K%(MC|p��S��&e�%��T1 ��,aݢ��O�Yjj}��dػ@!JAJ0#p;��vN����q+/�^[�5E$$��2e啩��f"��##�ʏ��db������Ϣܙ��=&>繁$I �ko����ߎ���!(�믿	��J�����[��W|@WB u5j&�7�FE(�2�p���a�Z�'GI�j8�҅,JR"��qZ�	����V�~n ��{$'�YTI8��:F��J�J(&��p�E�ZD���/�� ߢQ���џ�������a�ӳρN�BA]�:q4KU�H��bl�!���B 	y�e��&'Y4�Ժ�d�=*P(Q�<�O���y9��AQD�J�d��qi��~愤������ot��!�-��8R��S��������D�R�ҩԞ=�˥»�oV,;x�.�ĉwޮ6W�W	+�Kթ�� X���_�	��)��z��Q9g�ڽy��*'pM`+�嫀��%k�k :"�Q�_��R�/�)�����pK�:�*P�`K��7���r�D��}��D#!׮l������:x火�/oۺ����Z�d�RŲ'�V��'&VW���	�pa ^���d�U�
\+�s�g3I�`H�ID��G	%���/�w��v�6?Z�q8Pg4�L����Z���≒o����͡�\�x�~r��J��xta!��2��E�t�,d2\�N暰j��!Ō'GT��{B/�k��A���n����.&�NE�P4�b�xA/��
���:�1V�;R�I�5�r���-W:E@�~1WxU��􏎀 Pb�y&���5$�\� �UU�
��9i��,2Bc����`�w��S�>(��Q�|��;~�n7�/��%ᬜ�����b�"y�h&�Pt����K굹Ľ�M:�#l_��9E�u.E�B���\��M����뮻�z��׭�s����O���ܲo$lS����\Ν;�g�n�tHq��6�l.���w�K��x����={���
�|8V9�����]���<}�����z������ĩ;Hc{t�Z�����ᗪ^��R��SI�|����u���;*����]����%�P�B��jA=���`X�o��e�k�-��(����:�޵��~�,�����v�(�����._�+���	����K?��O������c�`��A�;��_��+�?�N������I���斧�~����ַ���zx�捕b1`���2L}Ǧa"68��ۻv�����CIAN	��9�ռ�.]�|� �cY�SUD���pg�ݷ/^�V��j�h����j䰜�Ř�{LG��Z&ʕk58G�jm޼�����1��C��7�/.��s����'�&�MӺ�}����y�ڙ3g��ȹ�g�����-��x&�T�����'���%e3��w����~8����㋃��#����#Ǐ��?�48x��G����=}��%�O,�L����/�p���@0��C��ڽ[��z=ٞ��X�.���+{�9؁���=�޻?g��6�#?|�J����r�X��Z�ѩ�E���=ǗTαAX���܌�~���nx���ЃX3�r���ٙٓ'O���[�y�}?�я/\��7�7�6n~�G
��ѣ?�>t��?b-P�{�=��/�:����oik۸��}�����vA(^ǎ��c����w������r�t���3�O?�wO}�ӏ,,.~�[߆J645�ؒv)�	�v��)�/F�v���T�U����#�VL
���R���)����I��x�w�%;��/n�O&� w�����>����~��v@&�7�D	����9s�R�b�p5o��f�Pػw/�e��7�H�D"7n��?��?{��۟�����|�s��B���+��șh�ٳg7o�����	^�~�z9;;�L��|�����7~���:�`+��
g�A0j�E�3���}����i�n�+�\���)�pjO�J�(;��?%�=5���A��d!�����-[���}��m7mݰq=�mjlnkk�x_~���|�3w�y�_��_]�����W^�+E(T�P�v��ڵ�P��>��C���PD�jb���\���<������k׮-..ʵfhe�\���t LX\?�@1��A�"M��\&�w;"K'Ҝ���H�򗿼���'5U�
�����W�qKU�wo����v�!�v�=�l۲}������7n@��m�A�
_y����o��ĉ���q���/����_��?�ln�{�����[��z�]w]z�g��>�O��ip����{�x������xv}}=�
Qv޼s�JO@5���;{�]�QVU������ya�HK8^�� ���N?��cpF�xTӸK͕m�4�&�硾;���������[o����wX&�5�_$e6L���(�c���[�n�C�x�I��?�$�����d�O��r�
�C���2 I��I�R6D�J>���=��7�	��裏NNN�.�_�˃so�
���e�tdQ�#3��ڶQ��!0�+_�J�T�#���^.�:�����_��j31�#)�s���s�|��E-��P~(
V�N�s�.v��O��f$v"��E�^�H ı	%�H�W<���p���O�Ē���
?��V#��,�H�°��E�z����q.[Ƹ���V&�_����?j��I��W�*�T�T*A��|<��L��L��s�bnn��[-�˔���D�)�J��́a�"?��]N��4W�dM��ħTtlS�s"�E�����O�x?��"�Ί��2�d0��l����`������_���D���jj)*7ܜ&΢I+�d_�ja��a����FGG�2K��k��o�hniinj^XZ��Tմ�W�A�h��GB�p�Z�7� ��؄�����֩����6�J�S�TWg��&����\>�-�����a�^�����"/����	'E���L��ӹ��H�������SO=���3y�E����=h�[��0�]����xTk%X����߿n &����]'�"����L��C���Ҋ�A�pS4����h�Hē�b!��ǣ�:�� pj��P[p0ljl���d"g���>�@'%]j��&�M�;&{=�27:������L��"�N��pDE��$j���0\KKc \�_����B�2:b&�g�[�֯��|��8�	�n���d{G[&��K�K/--�7�l6��M-�`��J)�L)j�2��ήr����U&�%á	.be�Q�� �P(�l�J$cx:H?�àF*�PW_'
�0�{e'�֮�+N+��PH�ke�bأ���/�I<j<�PZ�pi��@((g�s�7m@�466�Y��Z@�.k��Jޒ��XIl�تwZ�K)U��ugˡH��%b�����q!3#C���/�LۄV�*u����s���hhii�j�b	�NNNh��E[Z[N�>���Ю�5m�bl0��{)M�n�y{4�nI�Z��s���Ȣ�A-H��X;2|ݨS�x{S���Q�j�����PPw���������L6���~������O�)��V��������eDp׮]+qB���M�@��=Q[�2-�58H�}�<�rqk[��P� >^����S�\��'?�'�(�
S�~�%P�vB><���VhX~����*��m�榬���q�jX`���P��c�|~I��ΞB��җ���=}� Vuu����w�RT����Y�z�
o���������N�p�H�	�t��oQ��6�<��\/%G�Ŵ��!���k��T���G��
!"��80����G�5�pW�ٞ�����Ɲ;w^��'b�*����R��0�j�<=9~����3����_�-F��5]��VM�c1�Z^;(.��jҔ+�b�"yG���+_B��R)��<�W�PQ!��s��yS$U��!�;#.q�H��A�8$Oߛ�Ы)�([�Z/�:�((��C�2+�7�ߍ�H�=��p�?� ^���s�� ����m�7o�J'u��υ���o����@(�����Gn\������5�fk�[.���{���h��%9�a����R�qn�]V y�T*𞫌���n���̎�goe�'!�&ד��R�?���<̤��EՀ8*qd�k�V%�y�P ��O�H@;ۖ��x�������L0�tBzֺۢHH�I�@��������N��O=�������K}}��������ӧOG�q�r,��H����V�,�-5@��j �1.Jn�Iʜ���]urA���e�����1p�l%�(��Ԏ�J�_��I'>�Q�k�-��j% pEW�,�1��Hœ0� �,� M���D<��_���{���z*�k2���_H���ڛ���C����[�?��O��ٯ_+��_�_�r�h�v�.(�����r��.����#9�fwWw��x%�|�3EUR��Z���W��4VQ]�P)6����}��G$Bs�W.��t<�j�TCF�o[B�A⊈DW�4 $�����/>���u}�&��_|�j�����[�%(���_��Wa�/��r��h��pHt&����\fvv�T*�$�aóg��bNn��AX��D"����7�?Q۴T>W	���)�&�,F�8�����r|L�dv�O��%TLD�b4q�#�/"W�v�RL���J����uaVCScCC=>��x>�2�����;�S�t]]�.���I�u���������s���j��p�TH�4LJ�[j�X07� ���uq�a�N� �F{~	�i�C��tҲTߍ�G��a3�I0�"�(�oR�!�Ja�M}{�.���w8H19�[��E�Gt�>㝯�+@h�5��!��*��{	�$���V�X��^���!�p8��/�����o����&��)�X7��������6������^�$�Z�W���9Lw�Gw[m��!g2�HA��)�+�4O�X]L��1��}\��`{˕r(]WuuID��bl���{��wK;| ,Z�͓dq��a�vN���D��M�X{(�h�ey!4G�d����8���[�u�"���C^��F}��    IEND�B`�PK
     �;\;+z +z /   images/47e6ec23-9fd2-4f79-b93f-ab3ba2a25103.png�PNG

   IHDR  X  b   � ��   	pHYs  \F  \F�CA  ��IDATx��	�՝�/��QD���FPP@P6QP"r��~�F�$1f4'nY����d1�:�q4�&�!a4«�Qd���h��a���n��EU���[�����>/��vu��>���5�4h�����!�5���_?��G]h�7X��z��%�%����3"XB!�����B^�u�JcÆ��_��F�^�L]�:�r�-M�޽S��X�t<���d��+��Wu<�Fױ_�~�o��!��ױ�u����^mt�v#���ϼ?E����Y�~�y���M���s�e����[���v���o8Yw#�w����O<aD��v�I`�M�� �B	,!�B��H`	!�BFK!�"0XB!����B!���BQW_P�ʄCK!�(ɳ�>k���cXB!����B!���B!D`$��B!#�%�B	,!�B��H`	!�BFKb��5_Z͆��O?m�?[l���v�mM��:r=E2ox��V[me��K/�d֯__j0���3�$�qEK���o���>������ݻ��߿������[�[�g���c�X"B��R!��Ð�B!���B!D`$��B!#�%�B	,!�B��H`	!�BFK!�"0XB!����B!���B!D`$��B!#�%�B	,!�B��H`	!�BFK!�"0XB!����B!���B!D`$��B!#�%�B	,!�B��H`	!�BFK!�"0XB!����B!���B!D`$��B!#�%�B	,!�B��H`	!�BFK!�"0XB!����B!���B!D`$��B!#�%�B	,!�B��H`	!�BFK!�"0X��ٰa�y�嗍ho�|_}�U#��.$�D���;D{��y��'�B�	,!�B��H`	!�BFK!�"0XB!����B!���B!D`$��B!#�%�B	,!�B��H`	!�BFK!�"0XB!����B!���B!D`$��B!#�%ښ޽{�v�!�o^z�%���gn�W��ꫯf���[�>}���_�c�~��3��+��b^{���{��yܭ����w�߿�=�4���p-D;�'V�5LHLLY4z_ԃ~��e���(�h'$��B!#�%�B	,!�B��H`	!�BFK!�"0XB!����B!���B!D`$��B!#�%�B	,!�B��H`	!�BFK!�"0XB!����B!���B!D`$��B!#�%�B	,!�B��H`	!�BFK!�"0XB!����B!���B!D`$��B!#�%�B	,!�B��H`	!�BF��ݻ���W�^!��
Ͳ]��[om_B!��	,!�B��H`	!�BFK!�"0XB!����B!���B!D`$��B!#�%�B	,!�B��H`	!�BFK!�"0XB!����B!���B!D`$��B!#�%�B	,!�B��H`	!�BFK!�"0XB!
ӿ��;�N8��뮹>����s�-��´w0�y�{r��k���#�CK!Da���c_�2cƌ������[aS�q����f��Ѧw�޹>�7����l$��B��;��-���NS7^y��n�:3t�P����o��Jl��B��,]��̜9�8���{�1�j�*SGzzzr	��W_}�EK!Di^z�%��Ĝy晦W�^������k��f��ʕ+��ŋ̈́	���?l���#D	,!�A�"�_��_��NK��z���_l��>Sg.��r+ 'M���7���Zq)D	,!��X�|�OӧO7#G���y�?��fŊf���Vd��"kɒ%��#�4���z뭭�z��͢E��{�IH`	!��3�<c���J�"�ҮB���/ ˰�nMQ?$��BTƆL� q%� �%�B	,!�B��H`	!�BF��iT�F!D=x]يm�V�2y�ds�I'!����sϵ�E� �%�B	,!�B���=���?cD�y�G�2B!D8p�)���$#����i#Z�
bBQG���{����P!�"0XB!����B!���B!D`$��B!#�%�B	,!�B��H`	!�BFK!�"0X-�O�>f�-�4(U����^2/���B!���3���/��*�	���>���O>��v�̙c���j#�B8�O�nfΜYz;�\r�y�ᇍ�GK!�"0XB!����B!���B!D`$��B!#�%�B	,!�B��H`	!�BFK!�"0-X;<x��n����[om��j+��k��^x����5�>��y衇����7#�B��^�zY���7����?��y��`��mذ��^��FK=�<�@s��m��&�o8��~��}�<�Y�|��)�Bш�}��#F��Ç[#N�o�����B��[o-�7�.��bƍ�z�I�<w�m7�B].Z��<��sF!�"��C���c�������ꍦ	,v��C�V�2`��e�]LOO��ӟ�d�B!�{�6�&M2Æ+���z�)��1�cv�}� ��߿�9��c͍7�h��n#�BQ��X�p���{r}�)��v�,b�~�Y�~�,Y"<H.��(�<�W�$>�v��l��_�~f�-�������M��f[��	�l�-�5� �����Kv��߇]w��>gi�_l��_��Eh��ໟ~��G���;�lh���v������>k��+���k�#�i��춹�|�ms-���g1`��M�R{�����0���'��}�B�ƒ#�8���v?���?{�r�5r�H8��ν���F��,B'������3�QGefϞm��y#D��>��R۸��21��|�L�L�k֬�B 	��}��zꩧ���;ygq�AY�ໟ�?���.��eԨQV���.K`1�����G�!�B��{�=�,�$���r��_��s�]w��H�/����T��w�	U��n�)u�hW��yg�X��^{Y��������Go����P��"��CI}��	?)+�=���3�џ������\w�uF�:����Ꮓ�aҽ��RV�x`��E����n�QY��h"��ի�-eU����+欋Y�24����Aa&q#DX��i��i��=�ܳ���B=~�xo�Q����6�Q�j�ԩW�L�ra����'�}��ǬZ��<��F�P`m����4��{T\��#���/�����qb��g `��$�9�e���}�%K�4C��8q�Q�.��0��<�NÕ��4�+Ӹ�b۬R�������18b#���
+#�4���3lw�Z�L����Jr�N��,�e��
��h���c#��z�2�� ��d �Ԗ'~��L�>�̝;w3�9��ѣͼy���j�ȍ���������e˖%N�4'XI1�38�Z��8ӄ�	�4\f��â��:e��J�.�7%��D"�m���Z\�r�	�C����;��3��K�:�0�Bg	Ο;N�ˊ+�2���;�Ê7��(��g�
э��R�!	�Ҵi�r�DYz�����n�2��@�d>� �����JH�$PC�;�	k�³v�Z/k�7�^!`{��C4��H`e� �x�y�
I��V��8���I�*	�/Ci����`��A��V=!Dc�����z!E\m�6��h�T��b�N��7�7	��X��]7�{�a|�A�N<�����/���21+y����~r8�`+����;�e2bY+�<`W�X��lFfQ8�2�8z-Co[�* ��E]Y�K4VX�Ӻ�����s?vq��z��L`��Kb�}�-�],�̤z�Z�M`�F��*��A��/,���.4}4ވX����.1�ݬ�U�[+{\Q���$�V��dLycB�ER�:���;�U����5)�B��҄W��IXES�������g�ի��0(S*!JT<��T��ٞl��y�M�G��N!D1���/~Jo$	,�X%+-[T��������*i�f�BYb��9Z%"��x	\�!,��m
J�	!�6��e�F%+����P�oՊY�,�P�f��D"��V5-��G�T�oD��|�j=!�pU�XO���@� ���-�b�	T���c�m�i)7�ͥUz�g��,����}��m�!DX'��h��\�n�f�� W
��y�^b�&IAB�yՓ4��F䕍S"6��(����F#(��d}��cǎ�(j[���Ň��bS�X��<��h�z��ĉ�v��n�\�*J2$A`��#KR�֢S�Zo��
��W"�������x�8yI�M�
����v��2_!�`L,>��]�,&d�C���!�TZ1b�&�o�	����31��?������$i#o1b�f�`LHX�8紓��%`�溺k��E ��B��[dKr�ozӛ6�=���1�Fdq�6�r|�]�Y`m������q��Ro��˩,��U\��^?cƌ)�]��L��J�B��R�_@H�"L��3H Xx�bL�%D��U��� 0?X��q<3>5�HI��B�V9��e�,�*)���a��`B����e���J�S�&���yqͱb�Y܄��r��^Vo0n�-@}�Fe��JX��׋�{��JZe�"�B�!�'F��ڄ%��k�����A�?�����,]���݄��[VҠ�)E�B�$%l�hM6��n�Fb��ǹ#����9��r����L��=�,���*�I�8[X����/����-Q#��4�I��ޠ1{���WoT&�x���ݢE�̔)Sro�e�K��g�A�P��]�zW����7���E8�P�h��"�	gEa�f�@D�2n=3���!À�[�����C�D���%�3Z$��X��I�;�=^��"��lqΣ0�&^��o��6���.��Nr-�+2�Z�=���|��Ac�p?j�)��1c��9sf��\z饹@��A�e�2z�g�C�p��q�	,|���I�������� �����hG�\Cd?�ʘ͇���B`]��}vp�a�ndQC������#�4�^��Ij�ˑ�+^�5n	�zt�������t֥�Ço|`S�rE^�l�"�����!�p�/��`�9&D���`���K
c(�7Қ=�oDeX�r�IW&xR���s�`��R���2�[w!�@����&:`�u�H`!j�i�` "f��.�����K�=.=��*��]�^��:�g46�mK`	�%K���4���gҤI�Bm���I)X�|��R�E�>�xЭ� ^&�g��k�)m�B��J0��n��՟sT`E[��\o�ܰ� !��V��*5�k�P�2�@)�G�XΥZ�k)D;�Ho��%x�<�������F���1��T*� �'�i��p]��u�]ҟ	���$��k!:VP<nR�Φ*pM�A����O;�U�	,�]�@ܳ.���R�v$����F4��3�7����r�Ŏϛ7�̚5kce�,�f�]��M��$���g�@r�`��|��dڵ�XƐ�<z-��&D��Wo�3H��<T.�������2G}��=(�A|����T��D�S�!K3<�wgu�NT;	�hM+�P���UY�j�BoON\l^�"� ���W_mƏo`�f$P�����}f\�u��BL�5��
�|�c	���(!��Y�\)�<f����G]*�^�*�0Z�5i��.�8�<V(�fT,7�|�m8�A�(�F�,{��荢�)�&��	)YG8��Т�u�pʼ.�b�X����+e@�PT^Y&p�IE[��A�x��ƭX���Hj��C�V���>����&�;Mܺ�N�q�q%4�{��h�*HJM-�U��V1լ�Z����f^��@[�b��l��T��`@�?��xl_���[�!������j��R�J4�"-�O�\��߈^����y��� .���.�����<"���bE{2��9a���	a�Q��F��|��
����M�%���>��c_l�m3^9���m;:�#�X$��B4���3 �x.�z���b1޶D`9�R��301JL�N!�M��ި��`�m�>�I�X�r���#*�؏h��4\�*J�$���M������g	��SA_�q��7�0/-XIi�!DX��mě�j��^x���z�8��p?�F���!	s,έ�w BT"�\�wܞdR�&J��MZe�b%��8*�7����Uu��`����-�FP�mSZ&�8ܶń��>�o� "?yb4�P;�%D��JD{�*�%���u�zŤ��KB�	��>o;܇E2\���S��X�UB����Mp�C���.�7���y9�Bq�<;>�b� ���6�X��,v�5��#"���Y���+QQ_$��h��h���UT�GH��WQ=XB!����B!���B!D`$��B!T`�ACEң)�H�'i�4��BQE�#��^�2���!%�f�d�}�G�+�.��B�|(p���(پ�Q	]�/��:餓�Yg�e���[��|�s��e������VA����j�p�	�#�������g�m���}�v�a��b�.4��o�f�+!�B �N>�d�w��ְ�C��s�_��A�XPD�z뭶@"��Ҍ3̐!C�~�+�\����7�_��_�[��k�̙��9s6��b�|תU��Ŋ:65|�[�j�L�b��i���|B!D�C��o~󛶏(%r���[՝���Ç�C=Ԝy晶��'>���L`}���5��ַ6��O�S�����u���
���}�L�4Ɋ��:24V�`�_CWk�����D���_�����?7�￿m�H��:�˓}��Қ����B!�,_�|�К�4��Uft�EYq�l�2s�&j
����ޤ9{�	�4K��:6+�ȕ���7y�ds�ǚ���'��w�+�f�"r��=��c����{��C�ɵk����2K!���hP!I!@�����v�ڹ瞛��c>��6p�� �۔,B܇����C`!�����o~���o���߇�R!�����o^~��^�U�3A�� �#�<������+����E�YKf;��.�q��[%���QO3��zꩧ�#F�m-^��!��;!��5��k�L�,,R�s��ի��$a��)�w���,J4[����_s�)��`���r��,���i����~�Wژ02
�Bѝ��n�'��5��,X,^��^{٠�����C<!��9��o|�6N��ĉ�����y'���Z$����%�B�΄�uHs�����g�ߟ����V���T� !֥�}�c��=ѵz�j��;�#LOO��=��}��1�]w�-�����"|׻�e>����/���[qXB!Dw��
0�$A Ƕ�nkR8�,��`�C ���կ~՜~��	,�����%�.C�^�/(�K.��Z�(	A�嗾�%#�B��Õ�� �x�l�ϟo_b�C�+hJ�ҥK�O�&��I�T�y��ٸ-\�'��U����:,��Bѝ��z��'���CiX�<$MX�$=�h-+�'8h܂T~wAi��/��/.���o{��J�Sk��7�B��3m�43}���ۡ
@�zZ� -A�,Xд�`�SZ�W
V�X�z`�X�fͲ��)���=8`� +�(q3 �(8Zw0E:�o���B!������Ωe	�6k?���lҨQ�l�⶛!���1��C�c����7V%��h��*ـ�jH1D!RW������q<�@��/~�Zm�����zkkB�a�z��m�!�Bt/�ۼ�����'�رc�Q��Pd
b� ��jI��C�`�q4u�T��C��/��f͚5��w�3�8��?+�� 5�8�8���n0_��W�t�B!D{�r�Js�i���|�#��9-s�0�?���/��A�R��鎸	fG5�}��fݺu^ۡ1�M7�d�}�}������)��`xz$��?��Y�jU[7�B!Dxz�!+��*�G�'.T����+�@%�S�lSI,N�����eL�D�B�:�.2UӾQkB!�5EK!�"0XB!����B!�LK��(_O�+2)J�L�	x�>�hD����B!�y�H�^{�eu�6�lc�F�޽���EK�|�<��A��%�B^4w>|�-����oo:Ԗ`���m��f�
	!�B4C�:蠍m��8��������3�<cK>Qf
�Q���!C��q�ƥ
�$8Aԫ8��l��E�S�B!��<v�es衇�ڜy���GaA荢���	,�p(V�2�瞶NOO��Ym-��/|�]�VD���L�D(r�g�_%E�0�R@��W_�쳬Z��kNN3r>��<�_�~�ō��}?�>�j��O�
��]w���l�C���O=��u�Wѝ ���^ZFl����p�ܱө��7�������s�5�p�(���� �=]��}��7�P����|\�����h{���Y�1�&���~p�SR��,8����;�l�7�7����r��.�_&^���}��c��s�h�
�����>���!���e�3e�ӧ���F<#��z�j#�/��;����T�t��-]��!�KSH��0psД�Ǆ'�b��,�E\`!�ț�B�>a��=&��u�]���191�g�P`"�w�b&j�$�&��iR�+WU��$~|L`<��]w�e'�P��L�N�Fa�f�E|�0b��yK�<�f@q�����+��~yL�|��O�P�X�V��L���\��>�����~�� ��u!�M�\8�5�E��	1˱�9���q��B	wG�`���Ox.�+�1�x$��,"����96l�FQEK�^��G��-�E܆<�h�<�WS*2��rpИ�x�e�jo�8�!���������c��b�`�� ���I3z/!��YI3� F���%K6{�MX��p<X�L�~D����VB|ǃU���%�����a?;e�DΊ�ZM!`��'��$��@ �_���:�C6�\,<L�\����c�q�����y�����f���:A�}��s��:���k���Uק��a�����y�������{�0Z�xqfb����޸@a?g$�s���q���'�[o�u��I����j�i��v��κDE��أ���+c����P�*�]x+V���L�kԨQ��{����g``q��I�Pu�Qf���A3����z���?�}�&U�K������=�}Ť�9ۈ�HbE�6�G��p�9�n�Jq˖��{��q&P����������=��T�.2�0a��i���'�x�H I��?��t��m9q�1�Yu�����q�1�g�&�c<@�����q8��Iz߁�O��.���ɵAx&��N\q͗-[��X��Q�7�X���7ߜx�܏X<ݹ`�O�ֱ_ܫ�"��&+�,73�!˵B�qo��\��C����(a��x����}�9��x:Y����b� ����Y��!Ҿ�J��4X]q2<�0�181�1�30%M(� �b�%�,S����.k�fR���|aBd��0a��?OT`a�Ȃ����b���ILb-�HXRxv�65�J�(�8�\R�W�/��b�r�If��SN`!(�D��n1�9�����	5�� ���'�z��bl:��쿱a�J7%�9��V'�5b<�Vg�IW2�Ӊ,\��G�;�m�)*M`qn9��7���	��E�>ϊ�b��wk��q��q�11����&M����T`��x���b5u�����,�k��6�lΪ��6o �ho\p-�Wހ�0;WHR�K#B�#�t!X����xp�b�`�r۪*2*��D�s���8Hs)F_D`Aԥ�V�q���s�s�P`�CD3FbيZ��wg}�tM��r0p>A�oY�XN`9���.֎}����w�&�3Cx���zb޼y����TW>A�	,�W�&��oڴi�|������ܹs7S���\`�{p��/j!�I��N����(+�Ύ.F�bc��r�Jp�]�8�3v��4�aE]~΂i.E�����FD��f9uq�ܧY��('�E#0\�Q�N4����/���2��,��uD@r�fX뢸�S�-��hiqW�3f�ȵ0fa� �ꪫ���I!)q*{2�+�(�X��LR3LxI�:�ZMuL�MHL
+��x��po9������2� 7[V&\�2����}q.F�+o�����l�D�5EEa4��T�8!�+։<Ķ˾�Z�|��
B��q��AZy�4�.,�2X�R�h˳�ĕ8l��Y@8�	,:מs�v�B<�h&ܫ�$�(��x?&O�l�:I���Ϣ2���-	e��w!�
qk'�A�8�V��s��W�I�L��v;�(�\	�m}�zI\��˴;��#�ʜ��	�e� z?gճ�t�7��cs'��E` q�'�BE�+Z먨�s  �"
qC,d�\�K ��8ʢ���r)z�E**8x� ָK1*0�
,�7���DǸ��9����Źv�gU���B�k�fLď%Ų9� ��2c�hk֬	b].� ����{�-n�����~g���,�q�Ea��:_U��l7���C�3��:X1��<d�E�$J&`�b�`b��d�h1�"�kyrex��E�k��A�W�|��i�\c,g�+�@�NQ�A�e��<���f�w�&y�s��ʊ�����P_�xV������w+J��+�}�&��J)8��P��4zn��wѿ�^��6�\;D0�Ͼg�� cI�;W����=Eka���NN��#i�eĕ͒$�e�C%��)�B�`�	�<��'	��`SQo�P|V�I��-\��Nz���_щ��" ȸʊ9B��-o��~�³�v��9W����,���ri�̐IK� ���L��ha׬	6�,n��M�a�o���P��kQ�"2���m �\v]��ω��K�	,�F����X��11!B�(s��{wEC)��.R�#��0�0��la�:��yU�x!�6��(��v���/�$�(H��}�~0X�>*
��Z^΍�Ĉ��e�HA��z�M7�v�`-�<������������~��C-���;Q�P�gW�q�6���&�3�������I�ZR��g,A�#�"��A<&�}�D�h���r*�dΥ��<@��E����W�htٛ�5Yq����>p]�8�fE�]�mF?ù�h�3�y��+M�j_�Z��^I�����h�$����?O��m���>��R��Jk��-J����fgr��$��Hbq@�7XP�h��'Z���",��bt��B����eՋW�e~wH�x��H|�X�	;M��gV�=�%�(�IN�ǐ$��$*��Ⱂ܃'ȜK1o�+�o�������L�M�
��9:YD���Fq�E�����qU��Xěa�rb�}h{��E�Dm��$�D����FB*�JV�C�aJێL�"������U��hv#��]f[������x�w6�-d�L����A�����c�r9E�!j���i��]J��J
p���X�CԿB�G�.�2��7�p�f!�Ή�4��F����r�\����
��t�6�p��Wv+�oV$�xi��2�E(G�i��C����[R����խ���������&�jH$��GLt��F=֪������;q�:���ݎI0&b�q�B��q�2���v��4����}?:X�	؏�aq^�\~�w�r傳}⯲��X W\O�4�Pכ��k�Qq�(�ZW���-p��&�dm3D4���+�^$�N��0%�ȣ�I���m$ᓙYY!eR�=FL E����݉�i�?�����'���
�rX]��9�¤L
�s���%�e��NX�X��(ji��a1p�?,����"q�8pb�L�+b���;��9�[d���~���!��M���M�5�v��F���+3����(��W�	C�?!B�=�0��\>�Զ�,I����K��"P���h�'+�$������A�h�l(gA���ƊB����&MP�_��X�:SU�&ib�8/L�����.�dB�ѺO��M�#�4�𬻱������p�-q�!l Z�=�dX�#.F3�@`�`�8�%~������!�� �*涟t��l���/$�)�F�!ڝ{�}�k�%�ʉG�L[�:��ϳ����h6!�K���)}Q���ɘ���J�xbb��j.-��a��R����� e]V�]w��1Ԏ0��d�by�N�LX'�Q��Ƃ@qZg�
-��Q�aÔ�b�>���:'����8���M�9�{�ưp���p� c5A�-&�B�:q<�ob�8n��
֩h<�����E�Լ8Qq�CY+I��e�&m�'�+���k��|~��V�����E8E�*�M��х'��4�U��pClN�8�&A�]�X�ئ� ?m�Ȃ{֧�a��|Ե�����v�j�S�L)��_��׵m��bƅ+�!s|֬Y�٬ipoQ(i�{I��T&�P~����v�JLL�p��5�&��9�=^��e���">���(�fa��΋�	�	����}�aUGds�'V�쇫����"l��a��I�J� T�X�t�w5�w��7�5���p��\�]@�q�S.�q�p�#Dhى:���Lq�m�S+��L)��k�>���ٍƫb�O�F���s���9F�E�q#���~�v�=�l}�>K���Yj��kg��\�A�
�f�}��9�����1G}�wy�j�U��L+I��.�&I��Xٱ�b`n�R\�`Aj�'�6n#����I�I�	1��z�a厥+���`�Ǣ� Ľ��yX�G�8��ꊴb}q-���֓�5 �|'�Cg���(=*�DX]BT��rY���� t�P#+ ��}���5�I��~��#>Y~7�+��Yp�<���-� D���j_1~͙3�Z��3f0.�%�1��-�iT*�܀�V�����3�3Q����a�������
Q�������qq�D�,nrqV#&UW!��ł��h�&:V�|��H�+������m�Λ7o^��-[����3�b�� �-4���� �8;׀}��s�B�/0����+k��^�3��k�lK��ߺ����'mU��n1�a�te�D+�(o6��S���F�#�|=�E�	u��{�Q�/^l�M���>���ٳ����qY�ya��>f�X���y!��T`�vZ�/��9Q�+�:7�鄬�u��%D�WC�h�:�r��20���&�!�� y�o�k�g\A֬��E@Ȗq}�y��B	�WTK� �D�%�3����o\����{����T��b�auN��O�P�U&A�0
!�B`���;�yX�p��V.� w�9��B4_tA�*b'�B� ���IY�x!�򺥛"���k����+rX\�<T�&�B���EK+�'L�P��&�Cb��զa��[n�Ŧ8"�lO�0L�Fp+�^�(�B�,H,!{�2:v��r�1HУ�IRi_�*���C�"�
��]M#Ҡ9A�LJX	!����,�e���^$����r�t�@o��[�ㄣ%ˁ2$H=��7�P!�"D�2�53�f楥+���`�B!��DO�XB!���B!D`$��B!#�%�B	,!�B��H`	!�B&���`�C��I�._��5d���N;�rO=��m��Ɩ[ni�.��R�v!��3��sh}C�=
�S��_�,5`� [3=�[�!��:�ç?���~���\�o~���_��lذa����{���g���wڃ�B�QZ�|�[߲�r����ٜx≹������ok�B�Y�������:�L�<�̜9Ӝ��f͚5��}o�F��.��"��?��ꔦ,�O<aV�\�����p�΁�����}n��|�4�w��4͞=�v�F�Q�~Ĉ����X�����M>�=��C�A/X�`��sR�Bљ�u��~f�=�4���}Eq�p~��_�iӦ�1cƘSN9�\v�e���v�mg.��B+�0����X�����>��������|�[�j~�_�{�g�{C��⊝~�{޳�I��w�}c��9s��WD��������x�VM���X�n�B!��{��ꫯ.����~���O�܏e�����g���:���0�����g�69�3�M7�d�<�K�d�_�|y��jJ��UW]er�}��*1*��P�����O2�
qf�6if]F`	!�q���*"���������|�\p��J��������QGe������{�M�"�u���»�s�ׅB!��Bb�Əo]�Č�w�y-\y\���,2���7�ǭQw�u��y�����4W\qE�B!�(�/~��x��۸n�v?��ϭ�����w��f��+�7yw!~D�u�Y�J��ڵk��ŋͲe�2S'�B!ʂ+�������G?jF�mB����o/��B��t�hm,�M���/Y�Ĝt�Ifذaf�ȑ���w��Z�����K�'�B!B�!ȁA��G-���X�s"�����o��<��������~g_;-ˀ��J�?��?�m���|��4B!��8p����?n�9x�N8��a#����s�9g��w�m7���ݜ|��6c���/����O>i�Y�BP�}��ֲ�5���9UT!��	Y�;찃�����`]�x�N=�T��Q*��§I$>�����p�-�IwD���o�)F\�B!D(�8���7�ycI�jN�2Ō7�
���G��ٔ,B�	"�H}$�=O1PDq[�Z�(u6���|��6�M!�pL�0��F�e޼y�Չ�t�ڣ%���/Xk����~�-@�C��`���?6�x�;�ԩSm���Tr_�~}�Uk�ĉ��9�~�:C����޻�v\�!��A\3ޟ�P�S�@���d@��Ex��O}�S��T�d��	,Z���W��V,\�П�/Z�ȶ�AD=��s��@\Q�Ν۱W!��� �Ӫ��}�0D�b�1��4��Q��5��N���z��~����H���~��F!�"4r�����j��������8im��X��y��g�I��X�2��vۍr뭷�O<�4��%�i��l�T�= �x��������M��B!ĕW^ic��B����g�W�N�Z� �̵��!���8W�@Wi�B�<�}1�t�R#�Bx�x��q��t��KS]�B!�݀�B!D`$��B!#�%�B��
�^�z�zW4�&s���Tl'-�,�^x���O��B!D`��k/�;��f�7z��m�/z!?�����g��}-X}���%�n��z�Ŀ�~���O*�������G�V���?!�B�F`��g�}�Ad��'A�������m��U�V����ꏢ4]`2�6OLVIp���u�q�پ�T}�0�B�y��.�#�5�@�+*�cBo5�4M`a��@�Z�a�=�4�f�2===�f	!�b3�x�a��>}����c�=���\�re��7E`q��s��}�݃l������]�	O!�Ǝk{� nC�Zh�<.æ,Td(q��1�_�^�,!�BX�U(q��s�=gV�X����֨Q��e��n�m��'����N8�w�}6�0	D�QGe�A?���F!��	1Wt��E�;��T)x��lg2	�8�ClO��;Q*X�|����S����뮻n��O�0��]��,[�,��3�B�w�d	!������sEI�	&�D;�6
��D:2)�@`;F���4i������G�T*�P{�dH��ԩSS�wp�F�iEص�^�Xk��6;Ｓw�F!�Bt��ojq��n�m��M����K���:�����+XX��a�f�iӦ��瀧O�n�Ν��rDU�sE�	!���H���r5c�[d�\�����*1���'�d5
x�L`Q�=n�D��"��3Lx˗/��=���l���W^1B!��)�J�.�<�ʁ0�<y�5�$��K���s�6*X�ْ����w!1Y/���&�G�!�x��N��15r<e*�*�R!D�/^\z;uN$<xp��qR��(£+8�I��2��K/	��e�J�u�{�I��vX� ���2K!��s���WYHJ#�����J���r�Y�V�wF�D`aMJ���	�<PS+I`��K!�Btis?���mç�_%+�9	IqY!�/�B��!m����8k�薸�)��Q*X����P�/�sH!��G���HH�Q����_�������V�]ѝ�@�&�	,�x1X�c�~�a��ꫯ������ߊ��ޠ	��j+���4ƅ�߷�L����gR�)}! <�PN�ްr���ea�z饗��O��o�J�B��a�O*2J���⣾��$�*�ǩ,��~=IQ���3fL��)e���BA���
���g_��2�C�-v,���_�|�z�)�Z/U�^j�h�$|�Fe�$�V�^m8����w�uW�rd��m�(��lX��q3"�x��X�����Kt+!���O�8ԇ�VU�lB<ni+���2��ӄ9���o��Vs�M���m/>� Bi@Yֽ�b�
+^��v?e�+�^,���[�r	�
h��F&K�,��s�g shR6�M7�df͚e��<�p��ą����L`q!~��D�ݺu�� 8v�X��q��5�&�֬Yc�\!n�'�|RK����Vg#�x�y!��}�Y������y�L��'N�Xz;w�qGm�`ܸq���>������>z���4U����+΅Ϣ�2�K�.�e�j_aqaСOP�(��R�9	�V�]Q,���nkI"��wP�
�?��nDb7[�*D8\�QR�+*�ϙ3�L�2�a�;�q��L�3�~�R�� B�԰a��Ƿ�����]��N;m\y�����b{R�zJsѢEF!�,�ۀ8)��W��x�駭k�C�����8mڴ��Y�̞=���>��qY�m�bC�}��g�������˗{?��
,@�0������V�Ze_���4>���O!���� �7/.;�#BBt�(
��D.w	-!ʁ@�߈#�g<�ox��x}�Ʉ7�	G�\`!��͛g��|O1���I��;�4B�V��^�7;�c��א0���qM`q�3
!6+���7��<�',�p扡�\`�>Ls��h��ߵr�J#��7��{@�"ĮJz�`p�a�f0Fh�"��������\e��� ��dP� ��*oq�,�<�5�\c�@����>�vI��� �XT%e�9����b�7�J����E�q�X�Z�>d\$��} ��B�|�\���A*Zw��1Wx�jӋ0�[n�Ŧ8"�l��t��_�v�ZTQsp���eBL�b�q].?�����;z�!�Cha�jU����?b��6"?dS�"�v����XC��m��fǅ�4U`94�ϟoW���7��6��l7�!�Xy�{�H����� LTJ���4�̀�cTpaɮ���vwp!"����͆��T,�d
!����X�l��1j�m��X�K�6�'���z��UK�eH�z4P=o���:$���X&,�,�x18"�?\[��ye`baGL"��V�y�;9��-���F!򃈢^f�ff�,¼�T`%!S�Ղ5k1�$�*D��	�,�/b���Bha��B�;����B�"F� x�(�®BP
�mT�hS;�%����=L�d��
+Bw ֝V���UKG\����M����¢�1�]�Z�4��w_� ����H`	�% �?p�$�Ɛ]Cc�"2�5�'q]�	�Yx�WX�#e�;��s�Z�t$5���#	\G\��m(D=���K�\B<>�Yap;器]�[R`�@lQ*�A����5�`��	:X���u�dbJZYSL���] qCj'�
˖o�t,6��f�� ��!�ZX�ʤ`���v�v�F�����ː���_�^��)�������7�-��R[�4�� ����[�E�V�w�p6Ӳ�w:Ԋ�PnP!Dy$���`�25*���	�����*�px�>���LL��{�1��6+��%���0��R`�)C�`�P�!���N�WL/	JP���U'��(X��'��J\~E����S��Y�,�X"Kt+�/�ChT�E��xF�S��B�';���?��?��ɓ��8��H��BV�O*�	n�l5���Kj_�:,z��X���"�8��n�:�E���o;��3�e˖�K/��>�q�����SN9�\���.H��;��Ns��5k֘����^�S;�u��Zq��l� Z!�+9�Ti`&�=�u8d�κ��µ�H��UQ���5m�B֌1����ǲA�B�#+W����ujذa�裏6Gy�9묳lۜ(?����n�N�j�O�n�͛���<�|�D��~���ca�8�w�Y�h�@���M�� "HE��	�!-��u��;�C7	,BuȐ!v�ۯ�s���y��{ｱY�p���RvawC��E���.37�x�����}�+_1�ƍ3g�}�9��6�{���K.��|��5��z�-�<K���������w�5�J`q`���җ�d݄� ���/�ܺ#^W�@ �d����5���O�Q΂U11ZE�B���kV�{b��Rk��x�b�*���֎`�����o����m�wܺ�z�j��Ĝz�����5��I'�dݎ�V�2?��Os}omf9�s_��׬�B��KV��P�|�т� ���U��"K>�^U' �Y�׵�]K�9�Hr�;W!��3f�;�Ӝy�-\y��Z,V���;�����0B�b�B%�5��P�-�9^�ht\'����#K�U��:����۩:���A#L�n�8, �.��G?��9����b����_��;�R��k�����W�B�+o�b��Xp5)�����p�m���p�H��;,Yl�J�jb�tq%Bt�L=z�� �ٳgg.2���l�x.	����^�[>Rb��=Hp+:!D~����@�\�H��hS���@|衇r[�\6'��K9Pa�Ć��|��p���/l|���b���+�w��݆�w�p�u��Z*�H����?n&���ZbI
����a���~��v9yXMs}?��\��{a-�����d��RD��S� �����,D\I����~�����Õ��
,��8xLw�!Dc�d��d�b�Q����3��*��B=;�`���H��m��\�9����
~'1��S!YΕi`�B�:�.��"s�'�&���}�S����d`\%�C�G>����R��R:N�������!6�	3�c/l�I:jeI��u+����S%?o�1�_��A�Uu^Y��=e\�`!���mm�����6�;M,!�ƌ��$�#�82Q��䡥���oO��^�+�䐭S$��`�ゖ�F`�bغ�����L���d�@p��s?�8`���Xw����4�՝��8��C��q+��a,��-o�J( n��)�)����T�D9�[;�����f֬YV,M�0a��`<�Ї��s����@�_|���Ӷdɒ\��-X�B�A?����vt/B��M�4��v��!��}d��aboր���׃�B�`�w��u��A@R�m�B�<�d"���A�a�$�Ut6�C$����U;,���>�s�>��M��'?�I;}�߰�g�,�O>�ds������,B!D1X�PX4	&�E��yEm:�kX�ܫ�ٝ\'�<"ԕq��`�Y�L] !��_��W���ȑ#7�b��OV��P��}�{�򅻐�������>	,!ڔF֫vl�Y�� ���׀��l�V�?.C��$ @q��
Kq�X�U�]t<{xǰB�q�V`����~о���>19���g>��*$���OM��
,z�ze'��&�,��#�<b:���"��E�^YEU���Ȣ�U��K'��d�Y�Dv�i���B�
�X�e��������<������������*|�{�k�]����
��k�!D2Y͂YY���^W8.b�x!Xps�J]�u�
��������Y��]	.LwUK�;��kc�ҥK7�?-q'	���P[�%�H��$�^u�5��K�f�Z[X���Ŋ�ZW�ʊV�nDTd��.$����!�!�%D���RWZ�Z��@T(�7"B�sTg�"���Qy��։��u�p�B�B�0H`	�F0�fUm��ci���9�2�y�Q7ؿ�1s������1>�X��.D8$��h#p��Y.(�[�`m#���r�Dy�]r�#;hciv��G,E�iČ�IK
h5�'�7_��QÊ�ԡ���S�Q!��R����)�A�����&��,x�H�1�\��𜤑'���IW"�����ם�r/\]<�Xc�_l�� ^�SJ[�Ѣ���s�ǂ��D�4(�>0#D�%:�2�];+�Q��79��Pm�Z"��1b�-ߟ��ùAHkvEo��\�<!:	����""L�@��Pk�����Bl��y�����a��Z����B�,�G�1.�M�;c��z�N���=:� ��%��p��?ގ�e([#����L�f�O��	b�v�q��ޢE�ԨTtY�We-AX��`d}Oh\!Q^�"�7�TY>�sDI\���8�:eb��x�T�gLDd�S��z0	Ua����z�����n��cBo5�4M`��r�e�NҐ���===�f��­���*�qT���
R����I���劍�ʐ�BC��l>\�u�"�W�p�(^��~���aŒ����a�V*ۖ���k�f�\�2��"�8�c�9�d!`��A�x�jp,�܃i�C��p�Q��
YW)$>�&x1~���C��lTof �<��mȱr|X�|��G���ˊd�W,��Q(ڕ�cǚѣG��nC�Zh�<�������P���Ac�c�%Kt:<�i�^��Ї.-&���Ќ'�EC5+F����v��"͂�Cr�����'�����X��rJ\ŷ˳�b�
��T.�F�ew,V�.���%��N8�5-��I⨣�2�g϶���J�+op;V���޻�e| � �/�P��[e�ZX�ha��$��V=Ʒ���¢�YԜWվ���<�}�h'�� ��U���n��"ak6��ir�!�c���������>� '���8�"�0�їpٲe�;�l�w�d	щ ��30䩾Mus2exn:�k��#b��0 ��E��V�f!r���k�����ƒ7EA�"����	�LX�d�\�<L�0�&����.��4��N`{���M�4�>c>cL����
�b5u�Ԇ�DN�ȑ#��y��&��X����:�����_� �����&����X�8A�"�U�h&�#p�q�m�2��Y�d�X��Vؔ�)��L:X�]`lKy�^&�g��6ṟ7o^���B|��z�W&��^�'�oڴi���9��ӧ��s�n�D�"���4�;��k�g�U���(�Z������3�H ���� x,R��kX�b�e�(�wr�v!-�
�Ռ32��8<o����*q�%�:Y�ƕ��A���U��I�&��˗o�	��]�v!���ok��Nr���ٟU-b�h�<X\t��[c�s>`�c�^���28C��*)JK¥�G\9f�'O�F���[u=�L`afKb���/t�܅�dū=3�"�0�E�
�<�"�>`qJ�:1��XfX�d���t8�#�B�H�x��{���getV��yzN�f�1�h�>��V{����w�X�f�s���2M�y���\%}g�.�$�+�qV�I��n��?��Y�n�+�O��y�I��VRI7��f,;͛q�󉋎�+����B�?��2�Q�65��bX�j7�*Iiu���=�eĕ͒$�|ƀJ֤��**Mx�Z5I���΅H"��Xd���Q+�Vù�͆ی@�"Zg��hչ�"�"��r��խ��1�^UH!B�6Nb�*K�6|ZSU"�Ҿ��b@�ھ�D�=M�q�I�g��t�@ҵ	b��zLv׀P�V�,"+h��,��E\�X�$�D�I'C�N��ǈ��G�D`QC%��Cm�L�!!�HZ�+,/Y6�\�ٸs�� V)o�C��)�L|W+�����"�e\���&u�J��8�HH�Q��J3�����O!��U�u�ѳ���J2����A���D1BDq����x,�����
	�͊�KB�Qw��i���ۤxM~ߒ2d�u����H)��C@x��u +����&D�c7���&c2��VwY�6[d�$��| X���<�V�U�h�U�3�Tdz�~�inx�^��e�L��'0s̘1���2yҾS�N!��I�[a�ثb ��c�ɓe���E[�f��,\}\�s�}g�b���+O=��M:�CU��Ç��vZ2��ިL`1@%	�իW�8�p��]wݕ�^��h��zV�P^��ܫ�X���Ad1�!�����U���yޱ�I`����O�8���H�&d�&�|�*T&�8`�0�ab���m5��P(���I�6l�Lܥ��}�F���ٷ��h�b�x����.*���3��
p�0��ɢ*�
���wI+�����$DY��XI[�p&��t�Mf֬Y�cR�^�pa�%��o��L`��HNz�iZ�$0v�X��q��5�&�֬Yc�L��<*˜9s$�:�,���&�0`�!���b�j���O���Ɇĥ�k�ד������̙3Ko�K.	R�
Xp�ƍ��{<�===�裏��'��B\��_�q�^1��	,X�t�-3���[�b�Ms�OP�(��R�9	�V�]�,xf�\8Ym���V8����*D�/��%;i&��X�}�����,N+]�?J�?%�#Ĕ)S��KWi�t��_|�T`1 35lذ���m��y�k�u��؞T�ށ�\�h���ȚвV�,X�Y�s9��Eǋ�w/�$�lAd�����q��c3�P�ݧ�5�/ͭ��X��̀qh���fڴi��cݝ={�u�b�����%�T5,N�9���|�r�p�J ~�(�ַ�[�j�}̉r�v#��R<�i�Y`���[�ܵ�b2w/��Nm|�A��۞����L��\��_#�E�lSz!����{Ĉ���L�7���=ͽ�{_ޔ'�r��P�7o�2�	�͓��I��;�4BtY^Y�A�V(y��f:ςq kI�V�ʘ��̽��=�,i_w!׊��%&�xpS6���}�f	,�`�b<��Z����J\�y�M�p�a�#�,D�'H|�ʕ+��HV-��A��X�I����p^�\id���Bd��>n8`�#���fAF!.�	��#��]DU�"�0��>jԨ ��ⅸ���9�6���r�5�؃&����j��˺f3�,��Pu�˪Ҵ)���+P�Q����Ft�����;ȲU�}a|4h��8�1p��OS�W�.0�,Y��Z�'L�P��&[b��զa��[n�Ŧ8"��t�G���v���*R�v#��zЫ�24#Й�c�E��.�8�4�s�	�%	ǷI4�͊�����	���E?�,���W�(�%�"�v|�a4	z��v[�EeK������D�s_� ʠ�ʊTbN�����V��jk⠙}X�x�Z���U�XEG��|�&���Z�fX���WV��mV�co�E�����X½��|
[R����PX�<3��,Z�$A�TϛE(D'RW�E����!a<@d1 ��� Y�!5��)9�c�C�ǖ�U\�|����C0�!�%��p���7�0/�����"��y�b��0`a���yH8>,Z�f�}��mͧV��ϷM�w|Ƨ�TY�X�(�u2�Pm�^�SRC�/k'���qVY]3��� ���Cl1HeYժ��+QB�ՅL1$���-�_!=H����{���GK�|H`	QC�,���S��\�.���:"�H�F<'��լ�$�&ĒT����@� ̚�o�V,���%K`	�	,!jHQ��[6�
��fMBx�R�B�c=�b�Ӫl7�����J�1m���G��F�sIդ1	,!�!�%D)Z��G�J>Q��-\��'^Y�!D��F5���%�>�t;ē�6\.��s6���+*��VX
��H`	QC�,��A1�Q`����D�Q�{ʷ�x�!) ����
�V�k�C\����FَNLQ��Cp��j�,D>$���!e��#R��N &��<�(�BDo��Z�vma-�s�=mcXQ¾6#�AK�"��F`Y#��,+!:��,���6+Ҫ�sQW�X�\Py;X��8W1C-┊��M�5\�k8��8>�B�V�f�#�}V�"�B��E�L�ŴDa��qb��k�m��:���Yg���>M?�O!�������޴+x�,^X��vr@L�2|ӛ��t��E��{��I�$�Z���I��lP�S�z<c�k6l�Fk>:=�����_���#�<һ����ApjRc�5k�!��,׌O�����q�d����g^Ȭ�]��jf?C"��8����5kF�߁P�N�C1���y��X�P�/N|����6��9s̕W^i�V�L e5�~g��0���'2Ƙ�;�"%�@$f)��N���d5Sd!q����������
Z��V�� m��uk>����|���袋̤I��>���c�X�}����V�����O8�IIn-_�;֊VW9	�m������D5���g���q��s�=�W"׬���Uv�;�?�}�6��s�w�W����0�&h��	��+(��o;��c"6+�% �������ӿ+V3YcŒ��Zj#��;�8󖷼Ů�X��z��W��U��!:b�V�U$V��P;,=�V<�������4�4�Op-�A\�\/�UBAT�x��!)D��&�w��Z����{�5s��5˗//����8��)V{�Z�3Ƽ��4\p�[Bti�^�x�L�$����I�B�?C����<qYX�g���|�,0�XX]!Q!���8蠃��B���8s�L��_��|��_n�2d	�s�9fɒ%vB�4N ��g�m&N�h�����˒%���B�[m��w�A�d�СM/U�/�,2�@xr�U/��N�S�iw�-��J|XB�=�k_��-�@<4���x����O7'�p���_q����r��lٲM����@������ȑ#����6s�%�!��,��G`b�xwb�^&;��[�ɠ�,�kל��!��j��j]nB!�^��g?��&�c|���K�q瓟��9��S�O`��C���cֈ#��FVV^jFd މ"����k�&|-Y�1���c����X�@)±*��y���.D�B�^h-�<�>��X��L�%D��"#�H^�g��w!Ytͬ�,Y� �|*����F�2B�uC�4��%�£�W	V,	,!��eϋ�6�U��w���jW�l�����E:>+q�Y�`'	,~�@*R�Ku��d�c��F�ϱQX����E}�f�N�0��� ^�Kt6�aQp���EK'��
q�=yh��b���:�qP����-��b:�w����C%|	�����Q��;y�m:p�!�|��d�ٸldb�|.d 2�4��=�2\�&+�׿J>b���&ڏѣG�L����ή �")$�q��3ΰ�&!/�����:6�]v�����]w�e��L(�p�I'Y�Y���#D7�Ȏ����\��qbA�4kB������U�m2�|b9�bU"�KKt
�%��.�r���k�a��V����w����ou�.�%�<x��O��o}+���T`1�S����~�f�q�7�p����X�ɢ� �*�\I�+,X!`0a��%�@�N����w�O�%c�vb��!�+���U������+D�aA��x�߿��o�/X�h�&-r�G��?|��!��!+V�Ƚ/-X�,�L�bF�e�������(--��vXc�R+����X� �p�m������y">7@ձIX���QX\r�����yR/T�	���y晙���w�y6yذa6F��߰�{�1��A�,Q�����&���xC�d{��d񽈍v[V ��V���fA�H`עJ��ueB�SWM��Bl�ҥKs}1�>M���r�%�Ȇ��I�6.���%�b�P&�~����,�����`���擽G`9�s[%,z"6�5�)3V,	,!�"�%D�!�,��$��fT�F�(!���V/,Au��B��B�q��T���zr�tY t�ꡅB����m � ���b��*�M������!"���J���Z6��]�	���H`�R����-�݈�m b%I`����$�3";w�:2�Z%�H��\���m���47q���4,�X˄ah����A!+K�Ԭ�pw���>d��
ѩ�,��	qõC�5��X(�A��7;p�81D�OYD��J'㝏�������|1�J`�Nk?m�{X<��b����5��ġ�-Xr4p>|x�iڕl��=�=��v�]	�m�0�'U]��%��`��Pz�����B�c�(>��k$Hy�"�U��a��{�p��*]y�v�����E	m�:�Ԯ.K�x�Ǐ����U�ly�2צ�!C��q���(8A���;�8�jMI�:�D�������69b�c Â�T��*�˧�)�k[��#�U�-;�/��nxv=�P;>恰
�bBo5�4M`a��@�Z����f�2===�f��7Q�ˊ�קpe� 
�<�,���W`q��6�q^ҼE$��?{g%Ey��7� � ;Ȏ,þ�� �,�d��5�37z͢11^s���s�1nI��jL4�BPdQ����#˰�l*��ߛSs�����^��9}f���j�����<QH0�}ذai�{�I�8q���Z�re��gD`q��Ǐ���	
><��y��
X�b Y�
Ѱc��op\D��e!w,�Q��OD�Xf?ß�ϼ����] �C�À�iC�Zh� ߏ�,TdX�ʁ�&�Ǫ^�,Q,$JY��b�iԞXQ�8�2��u�,��>���H�^s)� 'q%�"Wa����Rd&a��9���D0�©��D�I�N�6m�<	r23f�)//ψ۱ن���l:.��
��D��L�2Q��'b�g�� ����RҕQ����!��'�D��������f��͛�0�.r�n����D*�8i����s;�|n)V��[ꫪ�2˖-s��!]H���,!�N ^Yjt؞���75Y,�(F�Ǥ�Ui2X�E)���A�x�3��WX,%��b�VZZj��3 �.��4��Ca��X-�7t�P������u�$b5jԨ�'Q>�^�zY6c��:������k?�6B�;D:�F�PG�׭<W���,��QCˏ��d�9&*�
��|�H-����c:u��Y^�����w�	���3g�j
�Rz����=2�E�
+7�=:P-<n�83mڴZ�UI�&D1@:��,FcG}����|����{�k""�E�s���4�d��Н:���s�#2��e��X�N�0!й��!�l��ɮ�G�>ᓕ�|������d�	��U*��3Bx������%D!@:���[��_� �%uOԇP�w������8�D��ڵk�TD�(3H&\8���#��+��WB�3�������Ke��w}Ĉ6�㶍�o��Nd�0��0�Y��.�&�I,��Y[�l1B:����n�!�FG!�2�D#���ns�����t���$)�(!��'2D�y�˭�#V��4��>�2��0�����
�1t�����5��U�@�4X�[�~��k��ڰa�����(�t�+��(>�PQ��Ţ+7ݺD.��B1NN�*)M5� �Z`��S��	�d�='��x!�O8���/���~�q>�EXP����r@��	,�׌%�����?�A��xҸ	,��2���܄�i+�D^M� � ��6�;L�M:�||'��ϩ�CTǯ�y*�=oD-��y����� _=�D0
����f��.^��c%���za>�0Bۉ�/D1A�E��ř��RPU��°Jཱ/�.�"�HuF)��F���s�+���.|����׵??=G�ċT��c�D`Q������ñ�
�<^��訉
z1��2�(�B����7~n�n�$��#��$�{�J�����#���"J���=�R�,�A��������� A-�W$�(�#�'DY#�ɾ�0��QF����i٨P�
�t"X.�J�B�󃛗���A�������Y�i`��*+>����\��)��U���"��KND«��E�z-?�Q��]AP�����&�+��N-DE�����d�s^��M�Λ�:~!�.Bg(m<����/��:�4�^S�b�/{��T[�Bm<��Lƃ�C(]�۲�����t���W`���ѴQ�P��V&��@IIIZ�F���GoD&�AnkժU�{��)�{�]��U9:�o!�<Y�Vw@5P�R�~FI�5aAV��7Q����v��"�9��?U��(@��cBOuu�=/��g��%��4E&�8`�0�Ér����=(�2��B�Q�r���<52a�1��)xN(^�D��[KT���N\j���+����b�0:���Kv��?ǎB�}<0V:�HF��EnB}�Ϧd�1�!*��z�iΟ?ߔ����s�s��u]T��sm2"X�g��v����U���}��Y�^"j���&����|%��L�2ż��+F7�ʝ�A70%U�ՙ�	#�T^#��QG��D�X۶m3B��@��_��~~����kz.��0hРZ��"�g�6cǎ�]
��B\y-׬Y������K�Z�y��Ɗ+�@W�%��G)Ι3ǳ8�a�F�a���H*/��$R�n'�(��9�eגrA`	!j��y_�'1r�Ȥ�"t	�ʫ�����
,VӜȻu�溝�&������t.
�"�plO��@i.\��!�	]f|g��s���"���S1���NXB�&��/^lF���zyy��С�5>�.�Ir�$P�i�&;�.Q�eEE��r�H ~�%���*++�8`>(��^�T{$ĩ0"�T!]�n��#}�j�{��J�`]�C��4={�t����p��[�Z��(R����=s�L[d�UK�q��~�m#���a��^ŝ,|X�Ŷ�9�ҦRXQ�>�:	=!r�XtC{E�c	R�I���a�(v�8i���,C����+W!�;Nk>Ö��A�-��r�ީs�z�E*�o�.���%!҃�A
�{���>�x!��vQfD`���ӧۃ�-�BW�h���n!r	�o���n@0P�H�#B��DWTB���H��d�=qF���6B�"kɒ%�|VZZ����!5Wd�rf���-Zd[Z�����hT�WUU����&��xuϰ�a�ŝ|ψ0EŊ�o
B��\~K���!��>��:�V�|ce������@�{H����˓N�HDF�+�Y�f�U)"��q�A8�:���IW�ڵ�~@�LJX	�D���y	N<��r�Îb! ���í�:L�ԅ�>�X����utOqNMe���m�Y�%l���bx��b��#ڿ�~�78_�1="+�eH�zl�z�.B!Dr���cy��q?"�N4�
Ä�V*"�a�E�~"X~M
S%J��y��[~R�K�R�[E1����X�̠]�Aɪ�r#H��?|���B�%X�1"������ �R��������gAu�}T'yF$�r"�\\4�Y3QO��9�%����D�0��J:�$g�i��:/W�d �X~k,�Q`�Z���MP�������#�%D�A'."+Q�	b�H"�ZH҅A;�
ad�Jנ��Q����C��`aG謹��8�������u�B�GK�"у�!U�%���,Du�͛7�Ѥd��bvҁ����}1>+j�f���UD���&5Z�.o�֭WBD��E
�.�\��Db
���7�ÐnDj{���BM��0���^E5�}�X��d+��(�c茸R7��!�%D�\`I%y�E#���A�q�
���btq�G�2M���t#I�?����^�q:�[!Dr$��(rY����&#�u��Ȩ]Ӂh����҃���k߾}�4&�F��RW$�F�	,B�Ή�f i|�����WǙ�;w�l# ~�Ã��u>L4~#q~է��:07p�'�6Q�����M�\�s#�b ��{2�PjLy5�|O(� j���'gVII�����gz��u���������J#��.��_aѐ(zD��RN<X0�=z%jCON�~ˣX�T<�H��k֬Y�ǒ~D\�gP2�����z3j�([;�^x�<�䓵"�]�v5����i*�`���_��{�~L�\B�:����| �:4r!�?����D��"v7��m���n�0/��M#�e��o���(�8�1'�Ϡ�+8Wr1�SxO�jeD��9릛n�߭y��իW����.37�p�]��s�=�<���.�ù��%����޽{�����6w�qG`��u��x�������?���Q'�L�h���fCdQӓ,rCmR�.]l(��RX;v��=Da����+�W����8����S=D��H��Id��Ox� �ӧ�~ڼ�⋵�L�:�<��fҤI�瞳���=��B����m��f���js�7��⍣���k�+��P�am��<���cH�$��B�"D���Ʌ���Ds��S���<�!���4ç�}�	��oԈ+a�&�TLW����T@h��#89�TWW��Q�̘1ü��i�\v����]�����FƬO�>��D笿���V�$�s#�k�����K/�d�N��Q��*S��=Rg� ��,]G4�P<�T�HI���o�&WP��s�冸"������x�]��R`��q��[�9~.|f*f@�a&�Q����-M���B����
,�����$JWҵ�^k.��R�J�$M>�֊X"8t�IrN6^p�"��w��aXF���X� ��M����r���^�hq���UD�H�cg�����9�5)�MU�	Q� `������	)B�ӟ��5�*�X���GyĆ�M�շo_�aL�8�|����W#�V��Ir�O��Ӑ"u�(D����="eظqc-KT����ڌt@�8b�H�K��'w��g�>R�a��	QH �(G�����,�{�1�;&�u��~�����dU`90��Y���s`>��M9|��ߵ(��.�@��{2�����{������ z�{@�8�{�%��"�D$,
�H�"9������f

�θq��W\a�C��w���8��j������� ~ZƓU����_�rJ�;���{���D�~�_��@����ڵkm*����oNV���0�ĉ!��E�b��I#��}�O�<�'nV�,4�+�?��M!
�aÆYQ��
OM�3^��C8w����F����o�svAȪ��=��U��<H	`&�Q!rꢨ���.Ym�nD[(��a�Q��-�hY� �HYP����:2�VQ�,"��c��?���<ad�r�J�ϥ�y���V\�r�/}�<�쳁�ݳ*�h�&�Ή�k�(') !Dn�I��,B���c��C�Qg��0K��DYDP�>oΛ�I"1D�z�!!�$tɒ%)��j?�w�n'X���dA��q�;X�f�)�9�p?��$u$��4	�cK����E�4�~;����xnD�Z��|�U�����PNAj���\D�aLC��?_��h�{��mi��w�i�ϟ����}Јq�}�^y�+�(@{��Nن�=5	�XX%"cb�.S�L���قT�3��ZA"4,6�hq#�ET�2���ң�s6:�RU�g�+Y/�T��K�{y�<��S5&�zW��w�u��3gN���]�*) �H��EN|(YX�/~�� ���'Ջ/���r�-�1��k����<
I�"�����F��qN BF�|��Q�����)�Og�"�;�j*s
�(VH�#�8wPo�0���j=��lٲ�3M���pH	r��6�YȘ�s�z�g7�d]`q�����m��i���@��!�ӦM3B��aDמ#�HU�b�P��p^`�Id�H?3-B�5s,"X�rBc���*n*`"D�Y� C������ϟ"�NhU<�_�0�0(YX@��׾�53p�@ӳgO�$�@ޔU�"aEj��"��V�&����[�|BD5"ܜߝ!���#A�7����*��E�uԟ}�+!R�p��7'}Q�XH%b0� c1H�Eܖ-[lq|�89!���8�j��"��;�DgXe"��(�G�pbt����n�4�s�3��>����'D�mZ�tiJ�e��#+rF`	!�j�9�?B������F��Ät�*��U_%D�"�%������آ��\(�"݀�BX�j��"\$��9b�1u�7���( �$Ԁ9Q:�U�.D�!�%��9b�P_�Тv��x�D�NL�XA��VB�̑U��	�BW�6�à��"
Q)�$�NW��m���lP�>tr�(������3���=JN8���87ɧO�܇&�v��Y��b�sM-�n4����;������E�;������Nv�Νmm�˗/��:B���p'Z�#�8�8v�?�qR�M�9��%����bG�)�'D~A �C�v|F�n85�;v4�������fݺui٦d\`1,�v/a�����3�t��)L!Da��a	!�<��b]ك�}����m ��j`'c�#J�*Z�nm�����ٳ�B!D-�t�b���E���'Zo-F�%#�d�O�V�B�) z޼y6�'�BL��۷o(�"�Fڐ��#H�0#��r�	�Q��H�B!�\�%����I��+|?'r��l�X"Z�lYS�O'�S��pڴi��&t�5f�S^^n�f�BQ�PsE@'D�(zGw�7�N`f"o޼�vz1`� k�u�V_�'R�E!{���=�c���Ѽy�Z��}RoE�����N�v+A���5YB!�(>�$������6��{�!�h����
��:�y�СC��z?c�"X�=���D�F��t*=V�^���1c��V���MӦM�!�B�:u�a@@Q�d�d�M�3g�t��g����W�{d��Vn�=zt��~xܸqfڴi��#���+L!�ŅW���	&X�Q��:D�M�<ٵ���'|���G&�pgwe��"r�J�$^EEE�m^x��W�B!D�@IQ*7H�W�#Fؠ��6R�;w�L���a67�v���:�.�&�� �Y[�l1B!�(ڶm�z?)C��S�Bxt5Wn��5�EJ���@�������]_3�]?���\Hǒ߫�R!D�2k�,[��.Έ�\���+4����z�X"X�G�]���KxO-7��\��6c�Q�K!����0�氠���0�T���J�}�����za>���0�/�B�����d�q�}�[� ^�����
#�^��O:3��B�D�9QɄ�����?��a�_uHB!Dq�&�[�����@C�ɓ']�ϊM�G}d�(H���z#�vJ��޽�����B!���n&����2��p���=�Ⱥ���VeO�\�~�R�/�+{��B!D�p��;Z/\JJJ��7��?z#2��rX�V�2ݻwO�a�ڵ����w �B!
�����S]]m��R�&$��%��=�D&�8`�0����X7��`Y��g7Hƛ��g�uV�|�tl�lT�&�"f�qK�\�bf iB�n���盲�2{�#��Ν�Z�6�[2"X(��۷���6n�h���{|x��Q�W�6���W_}u���2e�y�W�B�@0cҤIi�穧�r5��h�A��چ�={�;vl��p/U�+���5k�X�dD&�`�ҥ�f���jŊ����vNP�*��9s<#4|[4"G!�(J��#7�+�!A��#G&-zG� ����h�C��!R�E�5Sݺus�Nn�(ۉ�4iҤ��
�Y���T3J3�1 B!��OH�-^�،=�u;E����C�v�uYN��5�6m26lpM:TTT�.G�T`��}��=Xee������s�۷�!��xA 1��gϞ��I%�n��>2l�?P��)r��P�9s�-2��*���BH���6B!�D�hk۶m�����r �E�0H��H����,�� �]+W�4B!��> �C�{�޽C�'/ĕ�̚CF`�0}�t{���:#;�.��B!����d��AXZZ���&�Cj�Ȗ��,B/P�-�-�-
��:�@�Q�_UUXE
!���X�n�5ń��5W~@cР�|�r��K��
,� g͚e�Ymڴ���9]�*lv��e? Z&%��B���,��Qh�ƍ[�U��H^����z���.YX(C��cՃv
!�B$�_f�gf�. dU`���P!�"�t�B�	,!�B�|GK!�"d$��B!BFK!�"d$��B!BFK!�"d�.�ʘ<�0B!�HF�F�L�֭��9���'3����h��>v�ƍ����U��k�믿��q�UW]e�B!��8���7�F�2�:u:eA�^x�<�䓵���n���/�~��;0��~<������~L��Ϟ=�s{�~���|��7�B!�u��17�t�P���3�W�6Ǐ7]�v5�]v���L����=��s�����̰a�������ŋ;}��8�	&�!C����z�\s�5�����OV�ɓ'͝w�麍�ׯ����}�ԩF!��ʉ�~�i��/��{�����O�I�&��{Ί)��K��?��v^a,�����3�<c:t�`��կ�_���O�k��3f�9��̚5kN� 
��[�����7V�Kh!��̝;׬X�"��0���}���q�md¸��ӧ�)��ԡ����`#^�{��~rV`}�s��?�L�b

�v��mo�,!�"�a,�)�!���:t��"Sy�CN
�V�Z��}�Z�1s�L#�B�*���߫��|?����q�I�E�j��^3G�5B!��r�m��(\EE�-~��vW\q��裏���?�5sN`�v�if�ĉ��BO
!�"Zƍg������s�Ѻ����&�կ~ev���usN`:�4k���ܹ�VE�B!�_JKKͽ��k�n��v�-�ѠA�qشiS[ ��?�9���9����~��|饗T�-�B���c���#��m�.C'bǎMyy�y��S~��X�G/������/!�B��P?������;�0K�,I��s�=�<�裦K�.�7�g?�YZ���X�au�`��g�Sp�����ɘ��,	!�(.���.���z��e~�a{}��~`�ϟ��9�!D�u���̚5��_�I��X�_~��YL��8�^}��i���W^1B!�#b^��bR)��4���{̊ʻ���&��"Ȉz1��+� g
bC4?jS!�οGyĜs�9f�ʕ�E��뮫�8&�,[����?��M����@�u��ٹ��!�r|�"g�S�>m�4�9!�B���?��Q�m����i+�bP�^=��o~��98�������6!�B� �ڵ��|��I�h�X(fG\%��?�~rF`UVV!�B�T`��ҥK?/�18~��%�BQ(H`	!�B���B!D�H`	!�B�LV��76mڴ�cr��������zR��m�6[�&�B�
�w�i׮���9�7N;�4�7��߿߼��;֏3�"����ٳ�)))�l�lذ��ٹsg;��J5VWW!�B�d��ļO�>ֈ����σ��W8`:�W�/��";�:��D,|@�a��}�v�p����B!
�f͚�!C��&M�z^�����m ��j`'c�0J�*Z�nm�����ٳ�B!D-�t�b��֐j2i'N��Z��	JF8~�xӪU�P��tpz޼y6�'�B4}��e_d�H�BsIfD`�"�W4!�cǎ)�%�B�
K\���ȑ#fŊ����b�"o,-[���짓�O>�N�6m�݄n �ƌc����ѣG�B!�j��$�HE����R�g��y�f�I�ŀ����֭[}��H������܎5F���km#�I��>�1���B�w�d	!��� ����
K���R�h�ccAt�HG�!6��q{��C��;v��x"X�=,� b5j�(��|X�z��"lƌ�~X�۷7M�65{��5B!�(.:u��iÀ���~��I��6AO̜9�US��գG_E�	,�WxX�Ao��с��9�q�ƙiӦ�R��Jr�0!�B^uWD�&L�`MF�B�A6y�d��#J���JV���=>�*"W��N"��UTT��v��3�<Ӝ8q�!��8���(���+�و#lP�m)ŝ;w&�Gd�0�]�vM�`HR�u���S�G�!��l�b�BQ�m���~R����
���
j��^3k����IӁ(ѱ��׻�f�	,������΄t,�u>!�(N,X�_�[�w�@vˍtĕ��M`y�f,�,�It��z�3��^A�S�M`9-��E��Bf-�#��B�x8`o�B׿�u=���J�}�����za>���0�/�B�����d�q�}�[� ^����b�`����:3��B�D�9QɄ�����?��a����]!��	��nݺ��u'O�t�?+6}���K� =��C�y�S��z%7�pB!�������2���|�/��?E��u��VeϬ�~����_#V�^�)�B��"~F��CYIIIZ�F���GoD&�AnkժU�{��)w#�]��U9"��`B!Da���x����WU�݄dܼ�W�'����x>��C�ˁ�{P��g����G���(�'���M����B!��/a{�*�$M��M8�|SVVf�:�@��:w�\��*�oɈL`��0�t�mܸѺ�8�����5�%�V�^m�&{_}��i�gʔ)�W^1B!�äI��-]�z�)W��\��`РA���EfϞmƎ[�.�D�ʫ�j͚5��?N���,]���̻)�+V�Ç�9Aɪ�Q�s�����Cآ9B!DQ��y_!	B�92i�;�q��LG����
,
Ϩ��֭��vr�D�����&M��xY�p��±=�jFi.\��!��8!m�x�b3z�h�������:�:�e9iC\�lڴ�lذ!a�MEE��r�H ~�����ÁUVV�p�|P��@=׾}��B!���z��麝T"����#Æ��MAʑ"X��3g�"3ꮒA��/��~�m#�BA�~���m۶I많ʁ�� �h�, �Gh�"�0�/r��w�\��!�B ����{�e�D�W~3kX�=�����AS��j�(V�]R�%�B"kɒ%�����4e�MR��\�-˙Y�^��-Zd[Z����@�Q�_UUXE
!���X�n�5ń��5W~@cР�|�r��K��
,� g͚e�Ymڴ���9]�*lv��e? Z&%��B���,��Qh�ƍ�s�=���H^����z���.YX(C��cՃv
!�B$�_f�gf�. dU`���P!�"�t�B�	,!�B�|GK!�"d$��B!BFK!�"d$��B!BFK!�"drJ`a8ʀF<)pQ��^6|����u̞=g�#GN3��֯��?�N��.���>�@!DqӨQ#Ӻukkb��(��~�C��S���q��4UrB`5k���s�=v|��������W���Ld��{�0Ӧ�gV��c>��}\Rݺ��!C�7��1��Ih	!����믿ތ5�t���mL�y�̓O>Y�����_��M�n�LII�i߾��������w����1Y�q9�>���С�Y�p�y��W�}_��W�UW]e�4���?5�p�9�\����M2�~�[��V�,ZT�\wݻ�{��G!�(L�:�t�MV@͛7Ϭ^��?~�t���\v�e�n0͛7��Xf������u>z���_�~��'��ꫯ��
�x�m��L�~��̟��gSVVf&O�lD������o��tN����i淿md���C�KR�
!�(\����O�_|��ݻ��mS�N5O<�4i�y������k��<y�<��#�4��}C�	%��u����}��|ꩧj�PŇ�o��o泟�l�
���j+$�}�ݴ��s�N����y�ŕ�?��������aÓ�G��F!Dr�.]j�oߞ�~�c�u�o��㏻n{��7�R�>}��"��x=�쳡���
�V�Z��-[�#G��
�E�Y�[�Uh�F1�޽��Yhl�v�y����ǧ�~���̽��1u��g%�a���[�P,N�N>�4�1�9dU`QH�v�rDw��/4g�y����)S�0��c��Y��5�_~�!�~@0��^UU���̪�jذ��y��a��D�ȍR��y癃���w�Y�.��ς�I������!�I�ƛ(\EE�-~�YXT�ñc�\�#��8��s�9�#����^]7��;v�y睳L�!�"�ƍ3W\q�����2��YX}��$�n�'u��5�ǎ���UW�!�%�"!�����{�v��~{F²*�P�p���n'ru����R�������b�B!
�z�!�;�j���}��
�w�y��lҤ����M�ڟ����S�'Q4G�Q(�B�ѯ_?+�Ȅ�q�fɒ%YX�M"��ܱc�)����o���[F�/���	��ߧB���W�^����?�������>�*�(b�5k��җ�d����lÖ��@���B墋.2W^ye���������S����i�"�}
!D�1q�D�^�.8�;�I�����Mtw�}��;wn��K֝��OcFb
[�iӦ�ګo|�v�9S��*�/Q��rZ{��u�L���\'�z�N����� �����5&S��ШQ#;�ׁ�+W�c!��\w�u�����e�N��NC�;w�?[�n}����.��yAL�~��̍7�ho|@w�ygA;�D�ڷ��l�rV(�4�}s�j܅B�@��ݻ��������X�=��Ӯ];s뭷��{ʔ)�%� !��/|��1´m�������s�H#���+��l�v�{ݺ����!�"���|��I�6:��W���3-^��^��E�O�nDaҮ�Gf��c����MyD����M
!��0��֩�v�Z69#�D�SVv������������_����?0B!D�#�%2u�7�x�~&��7]x晟���ö�J!��$�DFAd}��GL�~�������Z������#�B�WH`��ж�	s�̡C��U��={�0�{�9㌓�~���]��MI�qS��ꭄB�YX�j4n�شi��\p�ֻs0:)z��lW��m�l�(<�L]r�{F!�����;�Z/�;�s@o�!����~;a���á�^V�g={�4%%%�^�z��iذ����>X�Ub:�N�B!��>r0-�ӧ�5"u�,�ر�<x��UԺu����̸�b4f^^��> V��߾}�Y�pah
S!��G�f�̐!C�� 4h��>����v2&��q�D���zWgϞ�h�B!jѥK3l�0szc?Ȥ1�o-у����?޴j�*���}�����͛gCxB!�0p�@ӷo�P�E��!Q-4G��aF*2,q��A�ú^�,!�B�
K\���ȑ#fŊ����b�"o,-[���짓�O>�N�6m�݄n �ƌc����ѣG�B��=�t�t8���{��<������&DP��"��"Q��;��K��={��͛m'�04[�n��~"X�����s;�|͛7����'�V�������k�W<|i	�Q�%��G�~p;����'N�z,6=B��R��+,JKKm�]���E#���4P��6ؙ�:��ر��w2R���c���Q�Fynw���ի�a3f�p��j߾�iڴ�ٻw�B�| �ES��I8�(�ԩ���:p���@��'fΜ�)���ѣ������+<�� �7z��@���q�̴i�j��P��\`B!�(.�ꮈ\M�0������!�l��ɮ�G�>ᓕ,m���-���"r�J�$^EEE�m^x�9��3}���B��PRD��RzAĕ�lĈ6�㶍��Ν;�#2�E�͍�]��t���Ɋ/�D�!��l�b�BQ�m���~R����
���
j��^3k����IӁ(ѱ��׻�f�	,F M�2�:ӧ�%䷫A!D�@��8��۷��*d��HG\9�Y���k���"��֒KA���
�Zn�i��'_�V>�a!��=/�-]���k��i���D���k~��E"��^��o[r��B!D��u�2�8Ѿ�-���c�D`y���5�Ku���B!D���@D%R^D"�prX��r|B!Da�&�[�����@C����gŦᣏ>�v	�����!�vJ�P��FXN!���~7�Q��x����}����Od]���q��g�O�~�R�/�+{��B!D�p��;Z/\JJJ��7��?z#2��rX�V�2ݻwO�a�ڵ���%��,Z�ȼ��[F!D�o��cBOuu���J��������
������χ~h,X`�܃�e=C�� m�	��!]�M!��g�H�Э�p������̜u�Y���H��s��_��������ƍ�����}��Y�^"j���F!��,4��A�jmC�̞=ی;�V]��*ĕW�՚5k���t?�	,X�t���w��\�r�%��G)Ι3�3Dʇ�E#r�B���)?r���)#G�LZ�.A\y5ӑ�A��!R�E�5Sݺus�Nn�(ۙ]ؤI�/�>��
+��l�P�.4B!�(NH�-^�،=�u;E����C�v�uYN��5�6m26lpM:TTT�.G�T`��}��=Xee������s��$!�BD�q|={�t�N*��p���aC���� �H�,��̙3m�uW�RxMH���6B!�D��ׯoڶm���~��p�:�����}��(2c�"H}�ʕ+�B!��P�޻w�P�I�q�7����3L�>�4�h��ª���0��!���@d-Y��v�����Iꐚ+�e93�����8"�(lw�0t�F�~UUU`)�B��bݺu�R;�\��A�����m.U2*�h��5k��g@d�i���c�t"��eصk���h���B!�_�D�K�F�97nl�=��_,"Uxm�߿���x^�dE`9�)R�-T�E(�B�D~����A���U��Ʒ!��5��R�#r� ]���sK!r�Z�h�{�ЈCT>�Y��/V�9!� ��#ԩS�!r�|?����K1MV$���^�K�.�&�Xqꣅ$�r�!DnAM(b��wߵ�N$�WtIGU�!��S�NV`�<-� �%�>H$��sF�R�5"��D\���(�	,!����Ȓ�*L$�D�H`	!D bE��Ua�,��;J\���9�Ū�.LF�%��EY��x뭷$�
�� Q�F�u����Q\������RRRb�hjX�~}��YX�;w6cƌ1ݺu�7����n�0g!DNr��1�a�Y1���С��U������_oF�eӻ��y�̓O>�(���+�-��b��8l޼��{�v�_��c��ȑ#�X�ӱC��6���9^<\�9�������ݻ�~�D0�9b6m�$qU` ��\��*��x�M7Y5o�<�z�js��qӵkWs�e���M����=��S�W\q���;l7�>j�W0������?n��կ��۷z?YXp�`1�c�s�=g.��"#��Q^�h9p�o֬����>x_>��Y�t����*L$�
ʊ�~�i��/�d,S�N5O<�4i����H�z���D��3gδu�7�x�����?��ɺ��	^�,[�씉�x�|���5���ѣM�&M"}�+��bgeK�@⪰hذ�i߾��U�)0�&7�|�M{4h��ӧ�)�s	��7�x�F\9��0�\s�1b����u�%���1ꋢ����D⪸�1���h.^���s��Z�j�}L����믿���$�
���=�CX�tؐ�v��<��v������v{�B��֭[ML�8ѮXby��l�Z�XW�5跰��*.�>�l[SUUU�l���F!UWW[���K$�
N�\rI���C�=5lڶm��z��S�![��^��Æ��ƍ�5[K]��������xCG�������3��m��f���=ǽ��p���A��*p��B`щ5ݻw7ӧO}��kp�B,��<z�����jm'#د��� p��M˖-#�/]QӢE�;5���B�§����XQ*s���;w�z�P�%�_,?F��H`8Q	��J>0��N�Y=�E&޻B��B��C=dG\-_���q\cHR��s�k�V�ո�LuSE1�$������p�1c�ٷo����ҥ�)>Y����m۶ٛB"�M"�Ȃ` JӔ4SQ�U;����J��9p�@$��H4jQ�N!��#��MNg�l���իgǋYE����[�>��MS?������;����>���Ç����_>e��ݻw�� �U������ٱcG$���{�&�-[�!�(6z��ey�k�p�]w�9s�$}��ٳ���رcͯ�k;�a	6EXYY�Z����,�X�;8^H*��p�B#��?ŀ�(�y�5r{�T=e��#"�{'��%�K!��_5jd�Q|lw.��Bs�u��z�E�b8p=`��UW]e��1<���v���c�=��d]`5m������_�b��'O��J �`��vٸq�9q�D请gϞ��ARR�
,Ƒ�⁕�i�~��_�R�mC�^B�i�v�8'�/&�A`Du��$D��c%����y���OX@J�����o[s?݇X;x�'"�����o�9�c
=�|���ɔ9�<�E�`으  3�N.��L\B�|��K�!�q��&|�o~�;�/�!�LO��ݻk���G?��_D��s�\˜u�E!�>�O�t�}��z�j��  �ḏc�\,dHWO��k��u�%��M�Z|�R�s��	j?՚)�����1�#�*�B��V��`��?�')J�PP��X�df�C!�7����H`	!D�C���� ��o"�4g�iFÆS��Ʌ��}�5�0&&�ű�FK!r.�x����V#��7Du74�`}��[�K����y�lG6S0 nР���:t��ˣ4��E�dU`�G�ɠM�6��
�
�Z�2#]Cڈ� Fzd�9\!r"V�k��I-$L�z���%5��Ӿ�]�vVw�Eo8�.������iH��,VY={�4%%%�ҍ�ڟ�;w�+7N�P�ą��ٻw�k+�_�h��b�u�� �ӡCk\���0�;����
���֭K��<�뢋.���P�-��;+:LG�R�B�K��KG\9�:$ԩS'�R�� %:d��!�^�Fe6!� �F����	,�p(Q�thݺ�)++����B�)�Iz��� ��b���aÆ�F�T!�6q�D�^e�NP2"�8���ǛV�Z��?�
8h���	!D!�Ȓ�o��H�ռ����M߾}C�4҆D��A��X�ȰĕM�'E���eQy�!�(�Mg5/D>@�*,q�_�5�X���s"X�A�%�e˖5��tR;��M�6�nB7Ycƌ1���!�ǯ��%������T!��^E�BDi	�$�HE����R�g��y�f�I�ŀ����~�T`Q�޿��X3�a4o޼�6r��[ꫪ����^�.$|GM�"s�xr�{�����Xz�"����ߍpĢ2J��I`�B��^��+=JKKm�]���E#���,R���}�yC��u�nz$�Hj�9�C�jԨQ����z��eE،3\��ڷoo�6mj[����P9��8����H�&]� @���ye�(��Z@ ���_�~���M�3g�t��g����W�{d���+n�=zt�z xܸqfڴi��#���+L!�LP��lQ+D>�UwE�j	�d�/,d�'Ov-?"z�OV�EQd�4����3UD�R)�D�«������/�+�'N!��'2���(�%
J��R�AJ/��r@��1�uܶ�R��7�}���ѵkהցt!5Y8ǂ`Cda�W(pLg�uV�߆U�zّ
�v�Bdya�B��Pn�2ĝ=U(�GW�y��YX��� O�D����_���5E`!6մdV���G%:��x'BM�e��V�r2��E�u:r֮]kG����25��Z!������-q�fqX~|�"X\,݆�r��^A�S�M`��:rMl S�S��؎��@�ж���9��[�@�d*������(�%
���t�ڇ�q�,��C�뛓���\��`U�E��v�B�Q�n��kH�)�"�񺆄1���-��r��c�D`y���Z=y�'�]�sYl8��� �Ql�+D"h!?p�@d�?����H���k@2!�E$�k�CXc ����>/� 6��v�B$�I�&�%:��2�����Ap��{h�s+����4P�J�;������N�ݻw������'�ᐎ�(����{�����-Uh)�<C�\�k���(�oҝ^�>��3y!�.BVbnU���a�F���:�����(6R�v�B�����mhҁ��D!Cj��z��*PRR�־�,n���	,D���Z�j��޽{�]3�|�)G��)��g��Dt��
jF��a�}棤��"��ڏ	y<���֫*�� 7/���z&2��3�9�?��z���|u��i�0W}QSb����(��"UX|���	��e�P��I�R���af iB�k����MYYY`���s��u��b�-�	,�����]�v7n�!�����D��իM�PHb�!��(��"]Y���\��(��� E\ZZj#�t�b]@=4�T�z
x�9r��+|?� ������ٳ�رc}��!�W^�Wk֬�a�t(�ҥK=WP+V�0��s��U��0g��.A>�|qp/D���&:��x��;,Pq��GiD"�[���Za�y���ù�2���+�L�xĕ�[y>��y_qlS�L1#G�LZ�.A\y5�!N�/~��[H�5Sݺus�Nn�(ۙ]Ȋ��⢅�±=�<'���|��ņC��b:^�,�}q~�\���z��!Ū���S:P+|/^lF������rӡC���.�I�z�"���6$\���[��2�s�x����*++�8`>(�+����gr�B\p������9�\�aC�S�����?��X}����f�܄�A ��ٳ��v"{<��@���w��MAʑ"X��3g�"3?��A. ��~�m�/|��V���m���c���AP1bDM8�{1
B�
O�:՗��B�D�X�Ps�� ��D�H���H��4�9���h� ��Z�r�����r9�ҥ�kǮD��&�#����hӦ�)Y�d#���V�58Gԡ����0 ⅸ
Z��JH��O�n�B�Tga�@ۥ.B!Dm�P��.��ꫦ�@d-Y��v�A���&�Cj�Ȗ��,B/P�-�-�-R~S+4*����TL,���p"xQB��CA!D�n�:��ń�����Z4z˗/�i�J�����9k֬���S��t"�(޵k���h���B80#j�'��%���_�D�K�F�9�>�T���"REs@���#m�U��!E걅�A��B��!�9,��J%�$R�_f�gf�. �����sAú��y�X?:����2�v�B�܁�a����_eޤH��?��X�?�64ݺ47-�7Hk?���3��ږ�؎W!D�"��ǜv�g��}`v�6)�������˪b;^7.��Ӽy�;3łv�R�N�B��H`�9g�yzʢ����?j��xw��x[���C�/����&�1 �("�Y��Q�Qc�d><BQhH` ���|�x�&�6���5���������R�?�o|�F!�	��"븙��:�Iҙ��Q���b�"����Z��� �7�I�g����B�+Xęg�f*��i>�$��s�馴_s����]�?�Ʉ�+��B�?���u��֝�ڍ�;wڛB!D*ԫW���Ǐ���;v�QwLG�˗�+�0���7M����0`�?�����4B�ܢQ�Fva���"W P3a�ӵkWӭ[��iw�u��EӦM͏~�#s���r?���w�����^�.�>��ϛ������/��S���3�i|���͵�^�qB�Ψ	��1L��7��|�ߙ�B�07�t����Ǐ'�Yz��盧�z�f�V�^m^~�e��#F��Ç�_���V�0�/YX_����χz�����_����sw�W�x�!r�tB�Bx��O~bG�m޼�<���f�С	��A\�X��f���)S����۔����������/~�dU`�Z���^��}���V`1Z!�"k֬�� 83O?�t��9O>��X�_~�y�G��˪�"���jr��ś���={�!�B�0�|�E��w"^�?0LF������d�%�)B^�|��6,w�=�ԨC
ή��+���׿!�B�0�0��O>�����C��ZSh߾}~	�g�y�v"]}��f�ԩ6�GAZ�^�lt�{������2B!�aC]�ΝMϞ=Ͷm�N�֥K��u��o�*�e�� ��T%�:D��Ǿ���|��]�-��{�����&��w�=Ө!�%�	(��B>tA�?�UQQav��m�'-���~��qɺ�ɺ� �_�~�����g�m�f���o��fٲeFxs���f�������x���48��#�9�-;L����x�BD�/�`�;}��1�ӟ̒%Kl��D��'0�J��U��c�׿�u�S��|��ݻ���AL�6�:��������̿����j���6��!:b�7���/��B��[n������>�\_��¦VЌZV.��_�r�U,��Ϸ٩S's�9���߈SIE\9Ċ�|�؎W!D����o~co�\q�q,�Ղ��YXNe>��n �h�����b���]���������9��Y&�)��B�yb��z��m�5kfk�7l�h?YXΛ�袋L۶m�֭[O�>n�8+�(8;z����aˡ�,����x�Bd2gw�q���������BV֖-[�͐!C̣�>j����[��-r����{�9#��-JJJjڗ��EM���0kT!����/���^x���\A�PׂY�f�<��s���.�.��+죘$3w�\;6'(Y�"������"��s:������_[�/��-��E�T�u�]g.��R��9rDK9D�n���Z�_v�e�vb�Aطo�S��ɿ��/G� ��﷾�-�98�V���fѢEf߾}F�{�8q�F�R9�!D�)���Ç��oj�_�2�"�ň�خ]�R~/YX�LpB!�H~K�.�����3g��^rF`	!�CCH�F�j�M���L�@Z��	#"��j"�z�������T�o���">��"�8p��)nHKKKkj���[o�"�Hr'��6,���6�^�{��x��N��q��Vx�;��r	��H`e�؉�� �ZL�eo&����'�lᬂ��|�嗭10;M�41�w��� 쎈;]>vBd�����պ��k�5"sH`eV�s
�b��c�\L�[��9 �ܢbQ��Z���}EI*��*�� ��j����W2���cqoR��m۶����*t�+6��xEfa�5n)O!D~Bd�]�vVw�Go�v�iVop#u�1��0U�"�Hq����֫W��16�?�o�B�����˭}C>SȢ�Ml��
!���t����\�6łQ2t���<�:t�TVVZ��tlh2.��4h���r��I�&�y@xS��0�A!��Db�؎W!D�a� &�ԅ�A�f���6��H5��1�E�%j��[�6eee��>��Y�$:���b;^!DaA#ˋ/���8����ҥ������L�ĉ���ʕ+??#�?~�iժU(�;���Aϛ7φ��BA�F�o&��Φc�~����C�u�<G����`�����ޤ
4҆D��AR�X�ȰĕM�رc�de�T�F�o�	����s�̱�V-[��5�4��uC�)��.��ɚ5kjl��B�B��UX�*~�,JW�X��9�,��xc����T��IH(�N�6m�e���3f�)//7G�5�J>��t�F�o�`B<7?�~z~F���53~���:��+:� E�;�����J�9�	+�
Y�nݺ����T`���߿��v��0Xm�C�z+B}UUUfٲe�f��	�Q�����Cl��
!D��Q+.��R�o�>ۙ�%��ҀF3��M�65��s��5��j��d`��v�]��D�)l'����ڱc�/s�Hj/�u:"V�F������իW/+�f̘�z�k߾��O��:�����(��B�lù��)7#��}�]�����k&��G]'7'ғ�0��ˆE��:U�	z�Y�n��٣G_E�	,�Wԃ�Ao��с.��q�̴i�j)GT%9WX��ˢ#
�Ql�+��B�k2�|ƫ��Մ	�ɨ_��ɓ'��Q��OV�Tid�B[���\D�\�r1� �]QQQk3��<�Ls��	����Rl��
!�J��R�AJ/��r@��1�uܶ�RLV���"��F׮]S:X҅�d�=fD֖-[L!���\QRl�+�"ڶm�z?)C��S�Bxt5Wn��5�EJ���@�������]_�P :��B_l�+�"}�қ�+4����R�D`����֋�q���
�Zn+
�B^�~"P��?��"X^/̇�V����BQ<x]���<N�otK|A����D"��<8�58K���O��V!�BDC���LHy��b4G���ڿ��B!
4]�~�u'O�t�?+6�a�@Az����z�S�Z7�pB!�������2���|�/��7��x"�"d^�[�=�~����~Q�X�{��B!��3�'\JJJ��7��?z#2��rX�V�2ݻww�2��ڵk]�#��� F!�B\�1!�����zU��MH��K`yzb�L`q�a��YG,�n�A�����n�6�7BD��?)$�� U܍�������Eb�D��SO�������?3Ǆك���	ݺ	�ϟo����9)��;w�k��8�%#2���۾}�k�n�ƍ��8p�@����c֠��Z�z�Bd�w1�#2�$�Q�r��}6i��D	p%���mX�TkZd���f�ر��½@T!���֬Y��;2�K�.�'A7�+V�Ç�9Aɪ�Q�s�����C($w!�B��)?r�}ʔ)f�ȑI���%�+�f:���?D*�(<�f�[�n���m�b;�Y�:^V̥CX���fS��\�p�B!DqB�n���f��Ѯ�)J///7:t�w겜�!�j6m�d6l���t����]�����\�9������7�������z�}��!�B/$������u;�D��G��ʛ��#E.�J3gδEf~
R	������o�m���o߾5+@�L�̓|��"U�bկ_ߴm�6�c��Q9�"u��=r����Qd��E��.�
�=b�^ݽB�I�u(x�ݻw(�$ⅸ�YsȈ���O�n�B�Tga�@�%�[B!�� ��,Yb;��I�w��!5Wd�rf���E��G���n�n �HATUUV�B!�(.֭[gA1!%�C͕�4�-_��f�R%�ˁ6�Y�fY{DV�6ml!<&aN!�
[�]�v���I	+!�B�-A4��m��q������"R������������KV�ʐ"��B��]�B!��@D����0(YXn��H!�Q��0rN`	!�B�;XB!�!#�%�B2XB!�!#�%�B2XB!�!����(_y�1�b�.��52���us���R!��M�z���9��~���ԩcJJJ��h��ׯ_�ҘȈ�:��LYY��֭��ᦊ����G���'|��_l��nӬY���Y?��ϭ�B!�n��L�0�t����&M�����.;:W^y���[�T�͛7�{�׎�JFV�-̷��m��ɓ'�l�ѫW/��CY1��?��`ǎ�5�\c~�ӟZE��g!�& pbi޼�]аj#R|O�����f�޽v�"��ƀ�M7�dǸ����6*��+����q�v�ߣ�>j�W�����y����W��U�}��@�%#���/~�;�p۵�^[�$��%�x�����^z��G�
���b��ŋ�.ER�L�7n���\3����|�N�B�B��?��O�� ��yn�С	�C:��[o�#��`1��x�(����������KF־}��/��9�;w��=�<O�:��m��ͳb�.]L���� G!�fi�I��-'�%�����ѣG۬�o�Q#�Ȟ�51b�9���m��/9�E8p�@�s�ҥv�ϢE���<x��B!R��d�⡤�H?�!������o�
�:؟;w�t�^]]m�k��!2OϞ=m�6�}Q����_|�!D�����@o �ڷoh�9+�6lhz���4h`��g��ն�:ɯ����K/�|�#G$��9��7:����������]8v����G�ڟ�#";PJ�*��^!��F�
,�+���
�qB!�A�7��ǒ��Q�T���O�A�b�u�	���B��.� ��pt�_rV`mݺ��t\X�q�߶m��X`
#�0�<�,a*B�wj���x���$�i�&#��z�m۶I���K���k�ʕ�g߾}]��.�8!���ܨ��0��y�bM�>�NUhٲ�iܸ���AX8p��ر�
:!��E�z�-3|�pӯ_?���/���sW�޽k��=�X���ٳ�\t�E�=rٲe5۸{�u�#Dn@$1�-,\�0��jP�?f�����<��М���|?��,&�$)$����B�$��IT�c��1z+�B](͞=�:��;���׿>���\CR������Q^d���җ�TS;ҧO��{���뮳����Ϊ�������d�3m�:u2?��l�ғO>i�	!��L|����ze!�z��cÆv(p"񄸢>;�|���(8� F���x'�k8�2�Z�\ ���0�* 'v�"B��{������<��#v��X�2��~����#Aɘ���׾f�5kv�}��� J:~�i��M���o����g?���?�g�}���O2B%D�.��b����]��ĉVd1�-:�B���I���l�%�����Y���C"��� ��e�]fo@�;V`��?l�#�����5�3,����3˗/�^2&���?�#�*�k`���{�A\r�%VlQ�����;�!�����%k��ƍ���XO7~'rUh��B�H3A�D���A~�����F���̝;��TȘ�
Z�?���F!�+���R�`�[� 
��m޼�t��ѦWt��SZP����0NR�^�DA)̊5!�� R4�p�JÈ����%̛C\���W�&�B� P�@�h*5"�ٷo�M���
XB�V�Zٴ&������N�֭[!�AK!R��h
޷l�bDa��Q�:u<����CVń�>�i�Ɔe)"叚vX�AY!�E�8�p!D.���&��D��5��7�4C��i�'�R۵kW3m�ACz��8�u�BVŃ={�4%%%�~x� �D�I9�Q�P]]m�"`��x�ŋ[�FQ8жO3�СCO���w���g�c?�4/��h�Hl:d�����ifɸ�b̍�1�> X'M�d�<��
Ka
!D:`D�8/�;"
<��Æ˫�B��Ǐ_kd�3�ƙ#�*{��5� �
D!��z4h`gBo����_a8��U:PxXVVfg)�%��gf]2��pDd1�K��,Y��F6�2>�<�)fp�G�3�L�ĉm$s�ʕ��������	�p����S�"20-��/=z�0�0Iu���<D��1|�B�qMT�$e����K\9pЄ��+�%�B"Wa����2�gŊ����b=o,-[���짘�1�pڴi�Ѻ��3f�)//7G�5B!�(N��"��"Q��;��:����c�%%�T2Łf^�!R�E1]���=�c���Ѽy�Z��}RoE�����,[��u��B�w�d	!��� ����
Kf��h_�袑�NCl(lwkX�yt��ر��<�Hjϫ�ըQ��vf�a�����;p)ʳ
����QE�4�*��[�]c�%�XI������c��clQņEP@Di�c	1�������d�3�;���3���׵ׁ�{f۔�{����"��'���bv�+*��A!���C��6(���7o�w;h��رc5�Y�ZF)zOL`���*�xÆ�U���e�]̘1c(GT%9W�B!j���+"WÇ�&�Q!u� {��ˏ(}�'+_�{bw� �D��BZ'f��N���>|?h���G!��%ED�� �G\9f��A���H)���9����"�D�Νz�҅�da �����\0!�G�!D�h׮]��I��^(£+��
z��)� ȓ'n�c���|N	,!��q��,n��f{Î�� ��I�3ߋ�&0�x�F!J٭ �W4K��
{N/�,N�t�5x�ƍC�W8�	�J�%D5���ф��D����B� ®�D��%lQ��%"����H��/�B��!��g�q�m�[��a�����bE����~13��BQy$�9Q��T�,�.���T�s|B!Du�&hڴi��ǁ����>����4|��7����t��?����vʨ0)<�R	8!D~�Ym���)}��C��w�!�H��A&�4؄��F�m���'�.B��U�3�w��oň�}�s
!�C'c!�H�e˖��z~p�ڵkQ�F�Eo$&�AAkƌf���
�2�9s�#�+� F!�BT\�1!��x�b�UUh7!�0�����3����_m&L�`���e=C�� m�7B!Du��@҄A݄�.�1���!*��=����W܇x�Gb凹`P�n����_�~��ǇǬ�05s�L#�B�ڂ����C�<���f�wnP�
qV5{��Hu��	,�<y����6m�����m���G)�7.�K�A�B!Dm�ʏ���h�=z�2dHޢwt	�*���f=�KX�Q3եK����m��~f�����^V_~��V8���;P�'N4B!��MH۽���fذa��S�>j�(����:�e��!�j.\h�ϟ�tL�:5r9R�?-[�����>}��o��[��Z�t�B!D�@b,W����'��c���ȰELOyS�r��Bi�ر�Ȍ��|~�
!�7�x�!�B�j޼�i׮]�����#�E�0��{�H���Ȭ�y��wɇG!��A
�{��Y�m�B\Eͬ9�"� {��ܾi
�
��Um��n	!�BxAdM�4�v8�`�MR��\�-��,�0P/���mqDhQ��a���Y�f�V�B!��-�ΝkA1!%�C�U�4���6W(eX� �z�)kπ�j۶�-��$�u"��ex���Dˤ��B!��� ��X�6
ͱ�z뙵�^���H^�~���8�wŒ��r�)R����"B!��"
�L�gf�.¸�*����E(�BQq�!sK!��ґ�B!�(1XB!�%FK!���H`	!�B�	,!�B�����`�/����y�W�)v���B!��Z�k׮�Y�ff�ҥv����_��)���M�1�t����pS����;�4W_}u��6������Mǎ�	�G}dv�e#�B&Ŝp�	�C�z±d�s�%��^x���W�պuk�������l��q�ǚ:���'+} B!�Q���m��k/;��[n1����ԩ�9����_nN;�43q�Ē=_Y�����g$μy��a�f�;w�}���@��k�a|�A#�B�=zXqEY�Ga���?n�L�b���?�_��f���+�蜲,r���sO�5jT��7�tS#�B�!C�؟�>�h��rL�0��aQ�տ��R�.B!�BT5o������e�V`0@K!�"
+V��?�j�W_}u�s�-�(�sJ`	!���y��7���ݻ7���­����{�u�-�sJ`	!���y��'�1�clv�qG3nܸ���>�hӦM�o�J��B!����z��p�椓N2�]v�y�Wl�;6�^�"�/���d�)�%�B����n3o���9���M�>}L�~��{�g���J��W_Y��5T���B!DM��3��۪��j�Vp�Ygٟ�n�
	,!�B�L�q���C���F|�
	,!�B�,�'�`�̋/�h�ϟ_��M`���v�5������-�z�����޻w����-Z؟T������~�,^��!�B���_���5�9s��裏�Fmd��c�����|.%eXGy��p�W���[omo��E��8p�m��H;�S���`�	,!�B�AŬA?ӧO7���o���_��+��:��sCT��k�GyĶR���B!��9r��t����l��|�����^��~����W6�ś��;�coB!�(�m��-�Ye�UlmR˗/���J�o�1�&M��r�"w!�Bԃ'�j�m�1'�xb�c�.U��*7XB!����o��+Q8XB!�%FK�
c��W7�{l��?��C���4m�����~���>��!���?��|���Kj�J9R�ZIU`�\o��L۶mmE?_"�u�%�R�r���R`��a��-~f̘QR�<G�v���o��BT\�����;�l����ZݨQ#�E�sA�$�5kf�y/k�����O���o�����*��ƍ[Q+���Z��Yw�u�ώ;��I�)^}�Uy^	ƽI�֭[!DmB���wn�bq��7��Z�
|�32�b�-̀�}�s��-ʾ��k�-�4���VA�q��q�<q�Ē)L!�����;�!D%�����nk�_�X��:�v�����v�&���F�Zæ�njF��9B�HJQ�%��D�N�̠A�lZ�PȤ���f������_���eX���v�ʹiӦ$ۣȗ7��/��"xB)H��X!��_�~�c���iC�Zh�8�ò,Td�ĕ�7M�.&E��0fٲe�l�f!���\�J\��ˠ�iӦE���VϞ=��
���N�+V������Y;�5j����O��LRc�Ԏ-����"��"Q��;��.|��Y�hQ��]߾}m�[o���$*�(d�ӧO��X3�a0���O��͚5�L�2�
/?�	�Q�%D��J�Ϝ9sI�q2	z>��-�i��(W����v�s��&!:�i��=�㏿�n��lGe���B�a���C�������ѣ�aO>�d�V����@�%K�!���n��[�2o޼H}\�H���+W��'	,!DV�СC��:��͛���=1v��@M�V�n�"�'&�8�aa�aÆŪ����.f̘1."��ɹ"���H����ey.�b��bQ�oq$��"������í�hTH"�|����#J���ʗ1H��;{�
QE䪐�I�!��S�6�o�M61M�4�C*�ɣA�B�,@IQ� H��W�����mP'�>R���n�m$&��ѹs�ެ�t!5Y~�~"������aA�_�$����a�D:R!��8� H��^(£+�\�y��)� ȓQ*�cԛ=���v;`b�[.���	!��[A#�h� ���^XD���k�d��
�8�$����BQ݄]��@K�6���KD`�=1B)���/�B��!��g�q�m�[�ea�����
K]�*���bf	!���HRs ��	�0X_|�E�ߗj��!�B�h����a����A��>��o���v:Q������N��(��B!�RaX`�	�}3N&K��\��LFf>�D�ӻ�ĺ��TeϬ�޽{�]#V�a�)�B���:KZ�Qw��vZ`���ɓ�W\a� ����W��]��m4KQ�Fb$�f̘a��j��.�(0o-H9�CD�(�B����֘VN��|p�Ǆ���ŋ�WU�݄d��VX��Kb�7�f?_���0a�us���}����y�B�ڂt%i n�_|ь1¬��j�������?X�}��|$&�P~��N`�n���ͽ_�~��ǇǬ�05s�L#�B���ހ��J��'���߿���"O?���y�ԅ���B\��_͞=�|��wy���Vr�����M�f����9A���Q��ƍ��C���BQ<-Z���c�~�c��T�ʏ���pb=z�2dHޢwt	�*���f=�KX�Q3եK�����rq?��_�z�L��
�� �zJs�ĉF!��ì�J����/�l�x?E�F�2�o���C]�K�z@�������9�~�ԩ�ˑX��iٲe��������x�|PQ�Rϵt�R#�B����8��ݻ�O*��pWď��MqʑX��c��"3��A�-*��x�#�BA�y��]�vy���A���aG����#4G�Y)�/���z��׍B!��P�޳gϒl���*jf�Q��3<����MS�V��V�]R�%�B��5i�$�A8p���}7IRsE�,3��@����K���Ea{������f͊�"�BQ[̝;��bBJ`���(�1h�{��Wm�P�*��A>��S֞�նm[[�I��"DPa�@7-�VB!��
Z�hb	�(4�z�gg+:_,"U�N0c��sW,�,ʐ"uo�z�.B!�B�\ ����zf��"�K�+�8]�B!�����2'��B!*	,!�B�#�%�BQb$��B!J��B!D����A:t�`�Xc��~ǜ%|ǒ �7�܁�.�qa��i^�U[�l�I�R�k兩����B�����]�����52#�6�pCӦM{1[�t�u`M���V9����r��Z3�RÁ��_�ʚ�z���k����coo�=�4Æ[�w�2����n���#���^�y�s�M7!DmѩS';��uI���s��2*�;w��NI��.]��kt%�0�֭[�k�'�|b�z�-�=JI�'գ�:�:�l��+�Gt��[o5w�}��r�	�<90�B^j�C��������vvN$�n3�Q^���a�H�st��C�>G�__�p-��O~b��o?ӪU������f̘1�{���Œ��"ju�G����ʎ�A��޽{w3d�s�g�u�Y�\��F$i�$�󒀃�}��J���Ⱥ�k���{�m��0��~��g����m���Fmx"���.StZT$D���b���3��w�)z�X�:0��F���h�<�X�x�J�B�<ާO���#�
���	�?����c���?n���kH׮]Ͷ�nkN<�D{=<�s�~��G�\w�ufԨQ���'�����V���J��F����Z��e*�Ȁ��U�hѢ��:�R�؋e�60=z�����7�~��I>�����OA$e�\��+-F) �Q,;Ｓݶ�q.O<�D�� �~����?}����D}DwF�m*j����
+��L�b�=�\[K뇬ڡ�j�#��T�·�v[�}�\�w�}�ݺu��,���z����4���R�/��:�m,Z�(��ЬY�Pq%D���K���M���1 ���w�}m��Ug�yfh����7�h� 3E�A,_��
�,E��U]�D)��J�)E�� �y�T_���o��J��*�Z��M]���>��w���ϨJf9_��I)�"�,r�dɒD����H^��~X��R���_��^%@'�4�!,!jj�KAR5��z}��N ^]�p	e}�L
,"V�w�M�<��c��/�%��[���<7NnW#월��I5 $$ڍӢ\5wBd�R�w�����JA�^�J���J�D ���c9ɤ��ȌB����\~��F��g�}�A}�0I����;�\)
��.��x�~�xR��V"C^��pѴiӚ~�b�#�TK�sP�]IA&��u}>a��>���A�֠��:��L�]��>�V(�{��_�RS���~���J��u��������9�쳋��X{�9�S�	��SO-K����{�W��|��z�d]hT���C=d��K/���w�"|x*�`��r��G�ut�щ9���/��b��S#te!��s�5���[oX��WOP������o6؏�w0`@��"�� �����R�A�w��W�������[�\,��q�%tzE�����z����k�b���p��Rd]2%��nS�� '�tR�QBTI�J+���H���H��Θ1������Vjx}a�Y�e<(_@<��6xprs �KUҒ���N;������j��O�x�,C��_Оd������
J�D��%�?���\��P*������K!Du��*A:!���kKd�E&�혊v<���r���Į���������~��5dRMi��B�B���:+��7�l�ǩ,b/��B�8��̫��j���B��LKw%�b	!������w����ꌫ���,"+U�E�']�t�Q��c;7?X��K���a�6D'���oB���$e�ȑVXr�!�a������Qj��3Ɉ>�X$�B��*���qv�/��UW]%�%j�`� ;��D�B�}��g�&�ɋ��=!�	��6�	(F����J��7�P����
,�?�\�ڒ��uH��n��"{��ɓC���F7O)Zǅ"h	6%�{��?�BLaЌ+�+�T�w�N�B!�����3�>�h�ϓz��B!D�!�%D�@}��QN��\��}�<8V!�"�%D�@7m��\�WH`	!j 	,!*'LV]uU�erE��=(��RX����o۶�iٲ��.b #)�����7�Q!�".͚53�m���k����,X����pt�JA*��ݻ��]����Z+�1뮻��ٱcG[��\��"�B�ڂ@��onz��eZ�j��-Z؟��0�|���f���v:F���|�]`m�喦����*> �*��c��;'�La
!����p��8>L���:�v�����v�&���F�Z#8F�a�~�iE��yae�)����g�}X�O:!hu�lٲ��S��}~�xe�j�¶��U��D��1V�׿�e��v��v��HN�vp��6�ݴ�ꫛA��|�s�=g&M�dDeөS'�]3�L���n�:1!�KYo�?mڴ)��8Hx�X�ga��"�p�Ax|��'9���[T�<�y�X�7n\��#��|�r;I#��g͚e
I��4`6&%&��;����:��5���a�`��9*,H�☏�2,��BE�J\9xӄ�X]*�%��s'G�BA�"vԳ�M�Q(D�J%���e�6mڴ�����ٳ�}a��x��+�Y�rv�i�v'Νv�Ɍ5�$���D��H���A��
QJ��ʗf�E�;��EUq)���̢E�l�?��}�ڔ;s�������O�>��c���A���O���M��,�.$|GM�B�s�,ꕊ���"b��"7\�4iz��%KV�w�p]pA��3�j��W��@� �䪹�s8p�m��{�!�h����
��܂�c����QjX�=,� b5t����|X=z��"��'���j߾��`�쎗%x�,���Ū:t��=�?��O[D'�k!��-瓰"rQ8\��\��[H�+��b:w�l}�� 
Y�G�N$ž����/6_�u���M������:��N�����\r�%����fÀ���y��y��6AO�;6PS��t��-R�{b�/� �6,Vu?ox�]v1cƌi DP��\`Y�C1�s��By�L���K�q�i����]5��3�8Þ ���4_8��]�D8��uމ��sA�^�\����R
;o��������5� f��y\��K�ZW$auW,��k�#u� {��ˏ����/
���=hd���U!��3BxS�Nmp�&�lbO�Y8Y��~V,������{���=�P[���G�޽m���/7|p��r!jj.9aƁ��j��9��E(z\<԰|��7���V�����$�*($*J��R��W���<3x�`�	���"��HL`f��l!o�A��0.aL/�`"Ai��"r�	�����3r"�w�v���3g�9餓�Wg�����?�����B$�kӦM��Xţ�P�E�v�O�w�B�]��s�&��A���R�7o^�s�-�(������{���:�뮻����O9唕B����k�17�x�=J`	Q>X��**Bd"�A#�\��V�szID`M�x���5n*��@`��J��΋�������w|Y,h�w����B!��Oص�T��m#ʸ�DV��!�e�r�iøz��k���6Xw���B!Dt®�qf��6��_��{/���.�R͢
�N13�J9Y���Z�[�	&�����>
uo����n�w�?�~���^Q�|��
ŷ�BQ}$�9Q��T�\m]'��K��,���^z�%۹�׿���S���ȶ{>���փ�"xf��1��㏷�+�|�8t�ҥ�N�j��qj�>���BT\wiV���8�P����S�ip��(�Ǟ ��2*np��R	�b���`#T��9/0ՙg�iG�2Ĝx����/��m�����J��#qW��>k5r.���_�ـ�V[�dY��H�T"t����s��/����g�18.����_�gd�1�>TC��<#�� �Q>�0�Ѩ�� �X|$v�a^OP�=�~�}*#�6aϙ��x�A�}����[�����;�8sꩧZc4vd~�}��<HJM-�	A�c���*����N.X���M�u���?���|?��B:is]�8)�X]m���zV�9I`��&�]���2��}�}��T�Ե�����k�Q<�R�@@ŝb�If1  9��4H����� �G���~����:�� �5c���V[EV�~�
�8r�H{ā���~�����8#Ҵr��(�pb�e�+/���C'
��A''�0�Ņ�m������`ԇ�	&T�����?�ԁ("�[�����s��0ՃI,�*��0���w��\�p�Ǆ����&$�&��=^X�a����Z�䏛{\8й0A�0+_��6�>"���B����μC�m�u\��|���B���h�6Q.��zc#����i nBR�#F����8�=�����{�Gb�ZZ��ŗ�E.*|x��D�̙3M��ٞς�"���s�F>ɉ�R.�%D�@��]��@�\�"%�Ъ�h`V_7�4����C�<��ӶS?��0�
qV5{��H��D&O�l�ւ���M�f�)<�W�Rdx؅�!m� x_?��O�sl�p�z��gͭ����!�UyP{����){��0R�Y����e�ET\�QP3N�G��f����%���f:��KX�Q3�=@<D���"��AX�pdS�@ifq������~F��4ω��ӨC�.�t��_ly�#�K�Dj/����v�R�����`�<q�^�P��>z�����=�ܓ��H>���S�aϵJ��bj6�u�V�E���
���/�l�x?E�F��iZ�X9Ϲ��j�s�?~�}}�ԩ�#���� ~Z�l:��7Fq��j������6��^{����.J�8B�}�����y�g�s��Z�}���UI)�ͼB�����}��*�p5�1D�Q���w[,J�W\�����.&�tlQ������ڋ+n��\ ��׽{�������0���sk��%�MqʑX%�6)2�R�&��`ܖ�r�ӟ�Ԋ���Ǜ_������	KlX#G��
\uY��� J����ӬY�J�-j�	�B���0)C�|p�c�e�r���E2��8����Ð�#4G���y��we1�O�{�aÑ����#�%��h1�{�m����(?���!���[�a���c"Ֆ����+����S����u(x�ٳgI�I�q7�^���s���M�+��Z�.I�djɸ@c���<V�=RXqݛ������x�;ɻ�p��\�8),��/�]K:�a-��@��z/r��h��s~��K���4i�$��\�P�M��\�-��,�0�������	*��F�'�,{��1@Q<2��B�B:mJ	u=a�Ƀ�u�E��n9��=~���o�k����p���q��[zT��j4��EL�h策Dq�	Bd�����!"�53�ƠA��W_�t���J�4�SO=e/��,:�܅�]���r���D��
0gs_F.�� ��2O�:M�@��D�s���b�͖�R��
�+d�)�3!!��.�Y�����	��@B�q�����C�c!���Y�%���8�s�uQY"U\{��Fo8�{�	"�Blj:�uq��_����������!K�~���ʎK�!��_!�?N�l�E�^��VHh�4ԅ��_h����|ˍ���BLq���b�����,E�8�p��5qN��J�[��}�L�gf�.¸d����;�8H�ْ�s�=��|�VJ�!'�J,pw���B�����wCw9y��8���{���?��Ǳm"bXrŨ�a�B$��Zk��h�DGq�-%��s�!c��5�Ŏ0�G�V5p�7ځ�X/ѹ뮻B�#]�<��c1�i�`�dE��T��8�E@8��9.�ȶ9!n��F6�[))c!Dv��W� 8�p_>�o!�"�� x[]q�欳�2'�|�9���mq?���!PӀ]"�K �u�5ט���Ê��D�p?��"�j�eb��V�Մ{~"��8����������1΅�9v!�"	�����{m'!F�Dxv�u���!��n�J*Ƭ8�A�H�gP��>����4(x���>��w)E"g4G ��`B���Q�~?�ǈ�+��n��5�f-�c��v
�������R��J���\1Кh���a���sϭ$j*���j����7H�W`!�Pauqr�N�!���1f�/�T�U���u/�sO�W)D-�=>a����$�\Q:����  y�IDATp�Ė�{�wD��)<"Ma+n��+��D)�.XBTD�]4�&$���b޼yF�R �%"C$�(�(7�C�~P��(�W`�:,�-�{�F!�PNd!�8���ȕ�%޲ �]�(�X\�)Z�{�u�q��3�A$ú��≎�0q�)��3�P�ӡNdQ��k�>��^!DmCI�x�W�2%db(;�۔�w�}�Zwz=I]`�}��f���j`BG����t�U�0����9r�y��gM�@,qs����r�3�ʨ0�/���C��D+=D�8r!DVA >�t���t�����9�c5E<���.
l���ꪫ��Þ㒺��С��X1g��>�*�7��n���w��l����#��E3e��"�\4
�����ډ>��b��C�a�w�X�g��c�=�t��i��n��Г�B�e�w��7%*����<&bE�Zi�XL�?`� ӳgOs�e��`P\����:������~����;�'���>�Q�0~�������위X�����vbo����N('�>� �`M��JƏ���ҧCTS�LQ�(x�����E��,���`N�a��W�t�M�3�0�r�9�c*O`�7&�Ÿ��0�����
9lg����o���"��ȢK'��B����8��.t��k߾����f&��/�)V��;��T�`k\4�0}X8������ٳ�-�������\".��\PT�-��'.P'ҷD�(�x���Ǆ	f�c]z1,�*��N����8�5�3��uQ-R�"|/���/���0�ER���qEZ�s,C�a\�H[�?,]HB!:$��J"W��Ϫ��`.��6�O�9s�d~� �ש��������bVD��E�\����s�b��I!�I�\���|����( �(ԫ���8��{"[n�e촸(���"&��%3��3�첋�Pn��6A��U� p����N8�<�Aw�ĉ��_l[A����"��AΪ*H qB@���7$�x��m+*���'���� o��qE������|X��]�S���W������_7�稰s�UΧX���k������c�6��w�3?�p��eF`�ƘU�E�5Q����S����w�y֘�y�{�*!�۽{ws衇ڂ~f�.\�\q;b�QЁ�#�0&U���]����A]�.��=��������F���bہY@8��ɕϋ��yyO<�D�mq��_!ܹh��r"�ψ�(]��a�6:v��>��7�4X�¾�ą�Ԃ��^�(=�����/�Ĭ�CV#����LL (BY��{�Ȍ�B5:�o����o���zk+B�7Wip��okƍg����o��$.�\P{�1����>��3�}\41䌒�J'��N��"j��N�D�C�#����my������e��ͬ��i�#�iƣ��[\�	,/�tdE�Wǅ�����$��kj����J�9��;t�P�oΧ�{��)�SO=�.��k�Cf�
����z��Q���G[�RIPT��_��|�կ~*��l�^/��R+,�S�{���n3i�O��X��!�x/�\}�-B�����o��&X`�����W��Z+!D�p�M��ּ���V\1����w�+��I��@� �HT?������/�y�Q� X��R!eHA�K/�dE%�i���7:D���P7�\ ������|��
���`���T)�B���h7�|[�I-a�,W��v�,.�1-=zt�l< �G-�sw"�Bm�{���z��c�=쭐΅R�����r"0�0ߪ$
3�l��������M��>O�U����b���ʯ���<���	���܂џ���A%n�I�9�T`��F��Z��i�&�
,7�.�Esq1b���k��f*	��	�zk`}�Q�bN!y���V�l����sϵ���%�A�X880U����q��0�K�|n����V�[��`���+���OMZ�yu�֭�ľ`���F���9�)�w'��3g�4ϬĚE!��c�ep���(���X���J"�_Nh��F��:�^�̈����ۺV����*��C����1cl�P) S��w_;�����o����9j���S\u��Gj�S�o�"_Y�	a~�rHc%�X�H��
a��+������pR��=�Z���q�>��tI���s���+tJD��Ϭ;SJ�������\��8������Ul��] �#O=�T�c���=�@�p�%� g.2�9����*�� ���Aޒ
k�v�D:�=z�����T2݄��	,�ȴ���'#'X���5sCٻ��wR�+�
0���H�I�&����IlCju>(��8�½���^�à���5H�	0a0g���������kԠ���0���r�)~�뮻��?�X\o���YHI
�h�4��*����� �E+;O)�d����@r)!0�s���~��H�Q�A^��]g!����~�/fx�I�x�w�r�K`	!�&ȿ/�82/,ҽ�-8��z<�T�b�6�u,��?���y�'�|�1/�s�������/>gJyX��F�E�(`6�j�E�:u�T/�H�w�q��c���W�⏨�g��]e 8��"S��;�vw#Iqu�Q҈B�ځů3z�â�_���J�I���D�s\Hr+%��j��&utN�0��o�w�ъ�����֜�R�ڵ��y�7����	K��(.�'��d�S�m;Q(�U}b��v-���Ҹ�bL�w!3r�X�B����b���z뭷�9��G��� �� ��-:���m�
�D��?��9�#�N;�d;	�"�(nw�@M�(��I�N4��`�T�K������R+��
�S#W���BF�$�EM��O	#��"���?����Z!�,�#�-�x�=��=�q�F��ڌ�Ym5�]/�����}��S�Bw��ChԨ�Y���B�q�&��Ͼ4M�ެ����[����^�BT?X	A�s�\s���:�����à�ᢋ.�Fwi��ٺ�oV_�C��7F�:q��ӈ<�]��X��NXk-���W�EAg�F�X!�x��݆_|��y_ !�	���"���y۶mm��H��I��R�����޳E㕘g�"�9���s�����رcth��E��,�:�L�}[������F�4���6ib��o��n<�J���٦�I������b������;p��6��//��r�7��()�wJ*��}�(�k���C��/:���O?m[=��ۡ�t"�}2��bK��M7�dS��d�8�˺o�+��aT�w.a(u�3�XN(�j�)��>?O�q��0���BQp]�+�W�^�U�V��iѢ��I�c��6�4}�t3w�ܢ�d�.��H�Q����b6cd0	+��,�}1��/y�v�|�Dcx/8t3�9��#|V�E������SH�"�~����ܶy^_.���2!D���1�w�ߟ��G�@A��b;'�E�+<����˸5�w\�	q�.4�S6��ŏ7JԪ��0���P�E�-Zdo��1��ۛ�BGNԄE��[S��s�m#��������3L��k��!�B�ʂ2�8 ȸ�ᡇ2�>��*jf"���w���j҉\�����A����i�4s�r)wQ:�K�@���������g����� ��:�;��y:_���.z���ۻT��)ԺD�:]ƍW5��D��ׯ��z�K�-���j�9�dA�"�P��W�4!<B����1�R���i[2���2�M���w|�Q��y<iP��D��s�PiDQT+<���_�Q���߳��F���SH��f��b"	BD��U�ĕ��c�ss�����>��\0��U�s�tn��KA���(���F��\��
�Y��ym�Ǐ��8���GmMG�I�����0�_~yf���ݐ�s(����%��xr"�����r�&��D~�Z����؋��B�}Ȳ���(���l��AJx�j�}������)�D)�>}��ޏ5]t~��PoE�o֬Yv�_P��B�����@(���o7�ڵ��ү��:�%�A�8	�q;����[n��d�,B��gN���� 
�.J��s�̼��K���G����/!��׃\5Wd6��B��_2�袌�NC�a(lj4���df��ۉ
,�^Xz���СC�o���ˇ{��'S�۷����2���C��9�������v��g ��]��=�뮻��X�r���_���/Au+�T�|�C|7�?��<^�B���/��a-��ra1�o��+R7�]�.��qy���Qp��A ����)h�U��4�nݺE*zOL`���*�xB������.f̘1�#[r��,�J�5��g?�Q�=���OH��SNYij7��Y];Ｓ]Λ7�d�n\��0�!�����Ⱦ��+	Q֏;���C+]8�2�P����]q�`�)e#Q!� {��ˏ(}�'+�u/1��;{P�#��B
9HY	M�:��}��l�.DۈRyE�hF������C`�בu�����!��N�:�rԏ�� ������j͚B��@IQ� H��W�����mP'�>R��k|�	,�lAt�ܹ�7� ]HM�wd
p��b�kz��ec��+�����8��J�vB�"��.ℋ�I*���w�U
s=����6��;{!e�;{�1GW�)	z��VX��<i1�":��9� ����E�c�(��w#u�})�K^a�:=��iX!Dq��
�q�@�	�������
�(��BG?X	,u����aZ�C���_B+��t���7 ����I�TE���2	���*��mD����
{b>�R\�rm?+>��݋�ޝ|������B�w�{Z�|����ӂ�7����޷�����:ē6%�J�*���`B�� ��g�q�me��~�%��w����Rm?KN�Dَ8���?�p�U�s�ǰvx
�]��z(��;�������b���=y�+�E=�n`��_�f��B���1�w��B�*�|\�@؉��"�g�t�m�,vH;��6~�.�n|��a���IRs��!ٓD������~���/�B�ظC;K"(_$��&��}"�������tb.�cj=�E:���K��������_�w[s>[��0��G1w�ygQ����hTN� ���X�(h���a������T� @"�H	�J�߳�k��
E�A�J���"?�XH�w�yǊ�|����I����FE!�	�� �Q���5��4�X!m�AU�����ݻ��r2��>�9�B����~�=����D]�n`-C�'���23��K*��0��Cj�k׮Em�D����B	�3f���ڪ����9s��[E!�A�ϸ��ۯ�;2-�= ���u�딨�΂��f��
�&Dt�	��@���o��a~(,�0a�us�E�}����|4M:�A��k��4���c���gu���k�$ʆ[Տ?�vk�C8�u�b�vr	�C�YM2��5��'�r�����rt�L�T�������f�&��e�%��i���.jP�JY���ʏ���cdps�ׯ_����1�/LD͜9�d��W_mfϞm��^�c�߿��1���/6iB�3N�WF9x-ӎ�f�N �����s�m!�J!���w�F�T�ˢp��P!��� �ڊa�ȏځ�yqVŵ��=Db&O�ls�A�ZӦM�r���wy�.A>�,8�;���󪫮
��9眕�1���w����O�T<�4"T*d�R!��-\�Q�M��G�6C��[�.A\�5�q�D�D!Q�Ej���.]���*�(���_ɭr�P"���"R&N�h�+5҃��\_³�>�����|�ȑ�O�>��BQ<n�}���.�K�.5���}��Ͱa��';3j�([�@9��K�� P�p�B[���}�ԩ�ˑX��A<����M�>�ހ7�5}C=W�d��a�barZ�%���4��F#�9�	�q|ݻw��,��� "����P��)q��P;v�-2��*qRT��x��%�@�]�c\���-D���`!��uA���`�ƿA����p�[0�!Av�f~�N_~�� ��{��G�:*.�q�RX@���Ef��������_7Y�}�a�7�|s��Q�޿B�..qN�B�:�]��0��B;a����N�cǎ���,u��P�:���ٳ$�$ⅸ��U��D�?��}���كUm��neg�@�0��9I���\ďH�������>/��B�sG��?�3��ܑr�kcA��G�r�~8i�$�A8p���}79wPs����,�0�����KV�#�(l�:� ŉ�"˲0� O�m���֓E=q���g�v�RX��SKT".��\�)|��*DH(�:��p�"F���s�ZCPLH	�LQ>؇Y���Eu��U`9h�|ꩧ�="���.Q�Rk��,�5��H��xn��>��3�^{m޿��EN�|�I��Q�.*��a5JꤚR#iÂ҉,�\�k��k"�Gg�K��I%��PVCP�Bp��|O�֯V�D����YBsP�F-���"R��&�T�>�R,RX�!;��P=na���̮��j�<�H�%�t�M�s�;��9�3�����\�U���m[FƔ��="@����ˉ�,�go�,��p#� r��B���	X<��c�>�s�wљ���J���L�gf�.¸d�S���Q�_��W��.3���я~dS�(c�w�L8	��ѣ�k�&�x�l��LBB�\��Z��xbp���F�Pi��I�c�!Sf�x�5s�Z��먣�2g�u��
!4�����z�!���Ǜ"��C��4)]�E�"�� 䵩��5����elѢ������3��҅H��+٠�"�L�(�1A�j@�x�c�����f�b�� �C��c?�۷�&?��S��� #a�g���	�A X��G�X�����_h(�3�w�}�����`�7`��p���Q�H`e�<[l��� V� Ҍ���I��c���4Ɂm�K�!�)���Ç�N���m��&p$b{/�c0`@��"�����С����!�z��!DC$�2 κtROq��BQ�H`%�DUY=�Je�I���"ГO>�Z5�ʦ7I'w!rA��*Q	��b��i�'
S�m	!D%R��I;�φs��0¤}�+F���5	Yj	>��3�A���	��z�u�����I'�d�x�t�~��C��(5���?�<��[���W�û�g��eB���F~�硩��G5O<�B�r�5��Vj�5��(��u��VO,X��v�JY���;(��.���@�P7�x�{�gޕ�-��bk!�9�k��j}���cjF��,�V/��{���/���O�J�
S��;-���jz�pb�"n��r�B��/���D�b�ΝM�.]�Wri�v��N_!�D���y���K/��,^�8�k)k�����l���F(��_�����+f��~�
���k����q��ߤ G�i�G�9���qp_�h�B!D�����0��22]�1b�4h��Vz��mĝ!B�����_̡��r��몫��+(P�cƌ1���`�X�D��� ��#"u�w���Hܟ��'��Yџ}��WB!D	�R�L#���^q�f����7�'O��k�,`2dd��@QF���C&��G�m�=�X3d�ӬY3�㇜*����#��,�kf��?�I�eL����iB��}��1���%,Nt���,�̆m�;L!��gnq�&��9���7�1={���Z2)���L�2Ŧ�gr�Y^��~{[;�A�wXt@��EԲV�/j�y&�B!�̬M!��60o�ZT�*�N?����Y܂_x��#D�X�3	���ګ�qB!���,(dYV�E�>>Ot�Ӥ�����.:��)^�֭�I�M/�"�J���?n�uX�\rI�߻N����p��B!D�������6t�]w����,D��E�K��u�Yg�_|���b�=���/�hyj��Ƴ�>�YcNZ�w�i����TK!�H�����m����Ǖ��R����LD'N�h[)11�x�+��,Z%���:�.=����,�`,$_s��1B!jƦ5�7�n4G1	�7�:�BC�-5R� n���1"����o�l~������B�m�Z�C*�W�|�&�XD��cH*F�&L��a��n�\i���!�"Τ�������$&h�x��SZ��"�^QY-�)7͛7���S���C���E�l�æ�����E�{����B!D1����֯�j2d�J{K�Ⓔ��������O9��@�y_e5=(��L8�L�>��u@3�1��A���Q�2�0�0f�A)h~kй���>��KFj*���\|���!���+�V[me�z�)[U���/:섰�6���+�ĤI�C�����СC��~�;�;&���[o!�(o����E��#���bdG�+Rsg�i�ǋ�PE]��6��4^!0����<��A_�0J�ꫯ��o4���׿.Z\A��n9,�I�q�b�!E��|0���;�c4�*����B!D���vf��,��:"�.�9c�S����ɱ�&�؟�6�[���Ƈ�(���M�>}l���s� ~���H\`���:餓�Gx��?X8�bv��p�a�F!��禬�Ϯ��jo���WG8��Zk�N8!p�t[fN`QC��+��T ."�H�t6����3R��ځ�:!�B�6��x�9�{��q��BҨe)r'����O�GB!D.H�N�<9��$e�z�B!D�!�%�BQb$��B!J��(+;v4ݺu[�w��PtH�r�I#��.�i74M�c�Y�X�l��F���A������A��}/ӦM�f���6*��g�y�Q����jf�=�l�{��0DŴ��O?ͻ����n;ӦM���ƫM�2�����m��������q3/��B��<v��w7q���;�D���Xm۶�;?���|�)����{��`�Y��,9t�����sϙ�.�(���N�����+��a{�������f��;6�l3s�9��{+v�7"Q�e�X���<�븠#k̘1��.��B~�?��s͎;���#�8�/��v�����;�3�<�^c��v�iv��<Y��=�yX�C�f����}���t�UW�z��Π�O!�"�p�e�s׮]C[#9�����4�\���r`���;'�}���6�~��|���n��
� �����o��B��6}�t+��=a�b��j;��[o�5�=���p~��o?�}v_{��+��+D%�_���X悶�[�����M7i���^�Yg��Ŵk��,Z����c!������o��̌;��͋/���9��g�����?�a�+L(Y�q~�я~d������Z�
:�y�\�R~A�߈lC ��|�z�2�Z�
|b����u�,�+j!���<'��qAd�8+L�t��lp��[w�A�0��K�.��?�rEB�oȐ!�G_���gΜ9v*@��� c�z>���C`�(x衇��
ǹ�"E�����5~���KW�6dL	�Qko��1i�^�8p#���e�Ɯu�Y����y�'���#i���v��-��bS�<�UW]e#YA�r߾}��b��| �ޛ��1)�"������v�&���F�Q�a�M7�+
ZE����3g�U&)c"Zqf����9b�+���B$)�;7D���ܹ�MR_u�y煖��f����l�������>�h�]L������\p��馛�@��_����ST�:u����5*xdS�rૅ��KYo��n�����R�M�
�;pUd�MP����,j�t"�l�Bd�9y@#L�0!����}��g��f�A��~D�1�&�E�ە,�ʧ_�~f뭷.ɶX��6$��戓2,��BE�J\9xӄ�ȁ+�U��&z�L�.SX���$� �~A�j�7�u̽d<S���@���:�RL\����؁ Bиyo���W�$%��|�o��jD�8n�|E���<��W�: rU*q��.���E!q��
��W�O'!Q'�踢�0D�N;�d��QZ~Ev 'N-P�J�O~��|��Gm�E�_~y�}�#� �C�+�~7�!�|�r[�J������z�0X9+*&Dn�lS8_���ҋ+BΕ�w,Y��F�i�r��=��(��,�FGdj��Y���܎�@o ���;ވ���8�3K9
�
,
����z?i>��~�}RoE��9At����VD�u(��xܼp�����������]�ʏ_���x��֓��'��[�ps�P��ؠ�ϑk��j��ȏ�0�.B��D��J`!�,�~�n�c��u���Q�M�<��E�B�%W���D,y�D�ttb�@a{P�(G���Az�O������C�����â���O=�jKڈ��߻k����A���]waQK��"N<����؟(��~���!�b�+Dm��}���/�K#�("���.r7�|�������%�ŹܛV�k���?��=p��8���0 ��w�w.�&��ri
��0ˎR����"zE�z���;�S����9�_9�*ɹ"�De@q)�;�뮻ζkSlJ�����D��}��97:����@p�0P����O����8����-n� �ù�.WW�R7N��+q�C�BT6auWD��Yt�Cك>�Q���H����5/�0 ��\�:�0#�Ǩ?��S�e|���K��LJ�N�H�%	a�3f�Z0�!D�puV��8�����U��\8�w�a���P�Z��p	���6�lS���r��(U���+�T�:A��R$ˑ��a� ��(��:Hr��&#ظH2�JT&{�q���O�7�i�$.d,Gf!�(�{L>�ا�+���t��7�/�����s�1�!����;\�0�~�嗍�\0���a�hh£+�s+�s�&��A���R�7o^�sJ`U6x�z衶����(��aP�A!;��!L�+a^�`�(d6(�k����ǍWb�ꫯ����?�C^�N]q�vq�튿�鮻�)!��i诱��Ʊ�%��n��a��q�@�	�������"�ԕAQb���](A˵\��Gg��X�w�qvN��c�9<s�<����	���|�Gڂ�7�xÎ�`���V[�t3pB�� 
� �0h?�QZQi�jݬY�!
��C��+��Ҏ�a�Eg �$i��I"��u0��P�� M3�8.���I��
QE�="MT6a�~"P���(��XaȮT�U��l�ɏ�dX��8�¤I�nF� �Y��
W���k���A.X�����x��p+�\F�a9@ �Y9�Z�vQ
���Q6��Ba��U�,�]�
�I��v|���;�4 �2�K;�D3�EW>8W�X�6a��83�sm���O�~�%����8�/����9$�'�|#,�byO�:��@��gn�3������۰�lN��k��U8��=���F[<��C0y�jǃ����_on��k���a� ��s�%Í��'��HD`y'�G�}����;I�6�81�+M�ʂ�u1M(\Uε]Th���q �T���S�i ��]+��	�J�D!l�B��B!*��A&�Xv���F�mE�'�EH(7�ʞbb��
�f
��pB!DmA��Ó�@׮]��v�\�(z#1��
Xt~��U��'f�)G�W��B!����{!4D��Ph7!�0���?1��f��'L�PP$��}��a��4!�BT�֒&�&�ctĈf��V��M�������+�s�r���B����=]�$�Ǭ�0�Z��BQ;��B0��Z3ZL��u�a �Wa�W�g϶v>�HL`-���y_M�6������s��U��1���C���BQ��� �+Lf.��|E���UX3�z�($*�(<�f�K�.����$���8���뼬�)AX��dS�@iN�8�!��6!m�L�aÆ�OQ:S���\��5.4����9:i�ԩ�ˑX���y;lnol�����a>(nQ��k�ҥFd��>خ(��A�i��=��ӎ�H����۴�i��)7�9	��3o�X��ӳg�Ķ?v���Er ��Խ{���I%�n��>2l�(P��)q��Pb'�Ȍ��|�G@H0ʨ����L
N��v��"�I�?��H�I�㌯jѢ�If&��J1�Eă(��۵k���Q�D�H�qtO\`�>V*��b�"o��.�Y��R������(�6J5Z*I����4��}�B6���3�DC�>�)J*L�*��6�uدJ�$ⅸ��Ys�E`���M�6*t�ê��Kj���¢���Ap2"�g����� X�J`	Q= �&M�d;Y�� uH�ٲ��"��K/�d[Z�G]!!Шܟ5kVl)�H�\'V(&��%M�&����ܹs�!(�;Q�h�[���'��m�O=���g@d�m����	�.B����eR�J�ʂ�V�+�!D�AK�B,a��Xo��l����"R���~h���]����C�B����"Bd��;��R-��șs%k��F�ch�Q'�ɂ��/����0.�����"�E8I�va��K"����~<Ē��#;f.�p�HQ\��v!�X��}���+i�a���Vɼ�:�O<1�1�>\r�%e}]|&�_��JT�]�pW3I��2'�DncR��n��4hP��8i'%�.��Bӹs�QFҺ:a���C=伌92��%\`��E��c�-���UW]e�%���(��D8,����MS#tO>�d���oQ=H`	!%��j{~!Dm"�%���V�?��8��k���X5I�\o��V��on$�*���z�v<�w�˗/�6t_��VqT���u�I��}�#_|�Ŷ�&�9V10�8��*�5�V��=`q�� ��1��"I���'�!҆v紅�g�}f���%K���Z�Q�H`U��%�Da8j� ���dJ`�iӺuk���` t.!*�,t62V�n9Y!���,��O~���~�Ҷ:f�s�=��^,+*��H�R�������5}�W����*�a�z�\P"�X�d��㡇
5��ꫯ��>�\�I)��9�{�;%>D��F�Wf���W?�A����ѵkW���Aš�s��3}�t�lٲ�����(�4�$����O>x�|������K��U���|���qӵ�nk�5�_߬����٦��f�gݿ��y���3�!�Q!C�Ӏ�Є	B���z]~8i�E�8����b��`ݾ}�T��1ÌW�����N��1��Rc��o����k�m����4]o}�ֆ�=��.�͛77묳N��Kt���J�c��H13�D~���	,�i���
�f�L�b�=�\��G5x&��z��W(�����q��RS�E�P�u'�^�|<c�Y���L���u"j�N�*D3hX����������9f���e�	��4��e�o�ƮtҸ�pr����M��8FD%5j�T��d�ň�7��q\�������%u"p�k��Of�4��.���í6ؠ��d5mjh�a�
�m�����eu�[�x�i��Ʀu�f�=�z�[���4�Y?�k���Fjg�}���t�;H(@=��3C�q제Ҝ'&*V�4�.X`������7�Fu�ئ{�m�m�Ѭ���y��]݅���;�^6S�x�l0p�~�0�q�v��H�a��c��g�ubi�.�����g֬�8��$�i�w�}j�ϘiOz�Lzt�i�����M뺋&Q-Q{��7RX�쳏�y�wD�u""�1��Y���צ��[�2�Y�e�X�i��Z�e�ʗ[Ǻ����3/]r��0�Ǧà�m�Y���C�T���o���<m��9Ӵ��׬�Ͼ�I̋]㵛������>�M���G��K.6����l^�;FOɟ��HKo�"�H����7�(�	���1s�߬_'�6?�(�z��Eo�i�6f�c�5��m{��w�es癞d6c%-�e�Yw!$�VȞ��)W�=�A������a^�1ܺUK��ǘ�7ؠ���f��	'�63���w�e��`6m�������,���f|���P��ļ�{��ݺ�V��UJ\SӢsg��/~if��W�ҟ�1+���٢K���<����Y�z}rRO���i��?G=`���۬;h{�J�����{��6kof�~�y��k���o�i�T��7RX�AX������#�l����>;��";�X8{�Yx�=�ӠA�y�~�=W�5�4=����{�����5�O;ݴ���!
����3̛��o��4̬ݣgb�դY3����Jw��u�p���f��7�!��4�F*˵����P`ֹs��������'����w�ݦ�;�f��$����b:t�1u�n�-7�fg�m�+AC�Z�������g�첳Y�[�ğo�F��V�i~���f���N��2W9i�T�sK�{�7����SOٛ��{W�� �F�2z�*����i�̧�_g^��|����P���/7o<8�t8�,⪞��R�C3���Ҽ��f�A�6~Q���7RQ-�/���x�����<��F������x�Ϊ��u�ݮ�/��y�v�y�ҋ͂^[���.B��p��ܳf�u�1-�0��E]���먟��/�Լի��2�ԤH�4�Fja!���{b[?nܸL�����˖�Ə7=8И�\�Wo��t��>��{�5�{���#!D4������WL�Ï0?�d��F�V��n�ʹ{�1�v��B�OZz#5�u�]w��������Ӝv�i�ꫯ�������}��M�7L�ulԷ������)SL����"?x�ͫ��u0Ь��y�&;6�&�hޚ1�t��߈�$-�����q{�ȑ��r�!�_�~��6�g϶���J7�d��n��|(�&`�}cٴi�����R�Ya��v5�{�t�n;�	��P��\:���jq�������p�O�~)���.��Ï�-���mC����H����믛#�8~��f���~x�/�����2386+�i��t����	o��g���S�Z��j��Y���:�U�5τ�x�.]͊Q�̲ŋ͆��!���"��R:�����믿��8�(懷�z���y�5ӎ���MM�`�͌���K��V)G�Er��7R_r������n�������lZw���0 �C	�X��6��:4�q|~K�,1����g�v�:���haŻ�ֽ�[u�VK�ѬY3�A��=Ԙ�ǒ�EҖ�d�1�Q�ƦM�^�_Ӧ�V��fD�Rn����r���{��G5B����Ӻ�`��w1+Lvhյ����3�2B�p�����%f��ۘ�2T�A��f�믙�X5A��Ff�����/L�-��:e���l�M�'�k�j8�糏>2�Z�6+~�֐���ۛ�4B�	�
�p��on��j0���������i��ƙkv ŰF��� l�߱B@��1K!�w���e˖�Z�Ӻc�y���!c�F�u/iE�y���UD�ОTa|����7ް���-��bj����o�f˖&kP�F�����O%��J,\����ӧO7��7u��j)[3ѨQ#���oX$�wT��"�%*��|mVm��dV�5�4��w�"�o��ʬ�V6My����|[wK`�R�����D�f�mf�Yg��ͥ��Q�Fu�S�E����jF���u��H-D���cx��M�*���f��@w8�A�,v)�fn!���Jۧ��7i������t����'��a�-���l��v�r��W_5���I���0�}���ԓ����������k�a�_�¤3�*7+��;����6��B���ˬ����_��b�@J�2�bj~�.��t�b.6�a2�����Ç���'N4˗/7��X�eK���{�%Wy�}�/��j�{Y�^�$D���B`�'؆�m0�>�e���|���	�x�&tc@  �PE�K�޵UҪ ��宷��{g���~Ι�mvvwv�s�)��rm�0�'�VY��B������,��U���Q.���\�q�ֵkה�Ou�Ա3v�X���\�V:��4��β#Fd�8�^>s�L{��7���N������Y�SNɩ���]�9j-Z�6 ���c�Wbm��ȩ����J��[� ?h�L�*��9I���m��Ŷlٲ�_�Y	X
W_��]���G���{5+������Cn��cǎY�8^���gb,�P��B����T���+Wh�`'�����v����AӰ�承���)����~��ӧ��j?�z�4�����P��ѣ95��t�f�;v�H�Y��v��U������xC��3ƷpU۰aì�������&�i�zc��uQQ�۴X��te��}�vWG&ަ�
Y�{�=��s�G��W�z�ܼ���CZطz���կ����o��m���X.Ъ��k���[o3��7�1]�tq��{����r�*�޽�6m����ڿP{n���NF�K��~�x��k�S�}����M���Ol�1���n��uΙ3ǐ�z�i�����ȑ�rb��hU�}V}k��$J ��O�d>��00'�	�C��-����$C8y�Z��nha��W�o�uU7Ј����cv�����F$h�R8���X�݋�[$���	j�ɯ��ꫯ��F�_Ze�g�C~��K����v<o���A۵t����b��f��޽��jj��&�cx��m�e��m���q�0��B�!�sƀ\�z��bf
u�7�MzO$���_Bp,��;��R�ݯޮ�.��^z饘�QC�zB���O?�=��1�I{����~��Mv��W�䍼�B[��sVTݦ7e/��
;����:�n� ���*�p�iӦ�]r�%q�i���d%Z�X�R��X]u��Ҽ�t�N*UN�4�-��O󸴺�x�LA0�W���T_A޶�Z�j��c�̟o�]}�HM��^�>����}֬�s�Úr���m�u��M=T���q�zV����#�����1���"��lL`k���1?�B�2����lUUUu>�ঐ���3�ۀɓ�������,7�:غ�:U�����;g���}�;z��e����7Z�������X4��H��Ԥ�����AF?��V���c~~h�]����?l͚5��.VtL��WlѓOڨ+���,V��ھ�>�����@z\}��cx���ٰK�hG�x���o��?�sY9�b-��D��ǈ�����	X
A�cT�����Q�\��Վm"�e�66a�L[��k6�����c���¶�yݦ�|U������F]p�m�7��sNV�TV��ٶ�����q��/������j����	X��,w�+ �{��,���O8����W^��
�4��`)T��V7�o��7�d-S�K@|�zY�iSm��oؐ�/��8p�v����@�\N�x٢�+����m�?O0��k��fϧ�t��q��PuodO��=l�TC����}�4�	�;vX��56���r[� �Oa�~6���]��/4-U��ք��[�ؑ�[l�-��)q�!�N	p4A�"Q��'���VUc�O������66�k_�U��f-;��n��d<ܠ���۵h������^�����v�u�����CϞ�y�p_��#�煝.�~Æۄ��q!���6ƨ�>���ّ�s@�rZh�(t�T*A����`u��̼J�g"^AQV�iN��K/����m��7�p� +<�]��r���O��g��ּ����/wsE KEH'Μie�vٺ7߰nÆY���:�OT���.[f-NifӮ�2��yL���1v�PV�J�Lh�X*++~o`C�
R=c,�*�L��dqqq̯�>�����\���\c[8p�u����D{��z��u�y��tK�Un�aկ���ϵ6;���T}�N��+V^}����|]=Y�Aֶ��ER���:�qu+�>�TV��=z��K.q5���t�W9���7��s&�U&P�I$���+`�\����������u��ZJ	��|���Ŝ����(hM��������k��������{�4k��>�n�O���mѲ�u��ņ��`m���:Ff͚��������nst ��������-�x"�jTM�q�{_ak��5v����0+R�����(͑i]}�t���FL��3=��/�~��$�R{��Cپ�v
�S�P��v���jU���7��U����~f"�,m�\�N����]p�)?�J�/Z�(��ԍW��(�1r�HwK�٥^ܹ�C��64Nm�\��&�G��y�R�3�<c@���Ra�D[}��1������Z�ru�'h{�fϞmH�z�47;�Ũ�ƕW^������wމ94��d.hXeee�e˖�ݕ,X`ӦMK����i��x���/  �� ���SGY���_w{'���z�-ۻwo̯�^�:a�Z�a�ng�X���#�}��lݺ�%�x��w����  �,M?�U�J=�/����[0QobII�͛7/n�R'�ҥK���X�E?�䓸��4��n�#F�t�*a*���Jc��֭s*�H�� �h�@��G�#�=���ڲOU޽��^�iF]۸qc�+V/^���!���U��J�k��U����B-Z�y��x4���@  �Mi���6a��Qǎ7A]J5�p��]��&�$#���_��7ް3fX�N��_�+Yz"�#7�[�'UTT$����V۲CF���Fp45��������7َ�H�:tR���rT	���w]w�.��M��D,�.Vft� /����9G�:S�Nm�'+6|�����dm/B�Y���+�;v�5Os/(�P���, '�� �ǰ�>��CW�J�
ڦYlV�Es�R�-��={�&�O�<�M4K�E�+�%K��呩t����~{R����[m����h�o�ۤ��1�T��L��d��Fz6l�`�����}9���~�z7�J=Y�ƍK�p�z��S�9���KV�GsKTc����we4�����-���6�T���~=Az�pSnH�!���9]��Uv��nZ*
�^(�V�%���ѣ�����l)D��
�z��r��&	X�QJ��y��P鑓3  ��r�jj���*�:�*YM�bIe!  @:�
V��X   aG�  ��Iu��T�\��m��T���/�A	��Iv�U��Jk����T��ߏڌ�pG�)--��a�T�D�Q����[_%Zm4%�
�5��$�&o*={�t��B%�h#`!0�>���g�y�݀|���Z>{���
  �g�,�?�i�ƽ�¡�
w���v����l�(����jy���j�l
� ]��7X��k���w��/�����g?�y���~�UV�1c��ܹ��ׇb������j0鲤��^z�%7U^^n   Zr1odm����/�ٳg�2��8����_��_\:�����;n�gU`�6;�s�]��n5׬Y�  DW�䍬,��Ν;�m��f��������=���J����{��w��{�v�Wڔ)S  DW.卬��^{���o���=�\�Gh��d�~��.I����"Mc�Z��ꫯ  ��\�Y	Xǎ��z�~�ӟ�w���,:t��?�MT{�G�_�  @t�R�������/v�7�ԩS�m���_U�e��ծ�  @"��7��4����������ݥJ���y��{�4�6
   \r%od���y�lŊ�+N�s�΍{_ժ�   �ȅ���J���w�����w�RO�&�ŢBa�  HVS獬��K���=�8�W��^�y�}����}��1  �T4u�h��x�;�����ov��bY�|�{;n�8�*���   YM�7�$`�Y���̙c]t�]s�51�?x۶mֿ�ꪫ��'�l�1�5k��$6  -M�7�$`Ƀ>����x�n����
@�T��nW�bÆq�Z���e�]f����  ��Ty���֭[�x��b<o���+�u�M7�?���_���~�}o�-l���nu�����>0  �ښ*o4Y������rI�u��q��Ӎ7�U �\r��զn�E����  @}M�7X�Te�ݻw���޽{������8�~�[�7ް�c�ژ1c����-�ܵk�-Y�Ķo�n   �r1o�v���n���d��D4o�?�F�r��'� ^��4'A]艬[�����oaԭ[7>|x��i/35�aӻwo�޽{�����&�y.�M��7�t���k��օ�D�{�={��-Lڶmk�f�r�j���US�e�}�-�$��6��뮻,l����ۈ#�oժU����� $F���ݓ�I�G��0�.�Ʉ+	s-�d���r�K�.n8!L���I�y@v5o��&M��Vȩ�eȐ!ֳgϸ�/))�'�x�,�#T��k׮q��^�z�8qb���x{�!�44��׺��P綾^�f�S\\l�!#G�����[X$3o'j4��bt.����3M�Uw��j[�j�>'N��}��l�R˖-�[��z?�3ܥ��{L-��5���i�m>R�~�V2���F=�:��2��URQ��J�scm���4��S�籱s�����oqG��V�(����n��֘�Y�re('�̀����v�͘1#�����?���?���k�B+�� ^��VTT��>j���:�Gz��I���u�ģ�/�z#��?�p�e��w��ݘ��J�;�����/*�'O�+��2�����מ~�i�2�ϼFUsi�zߴ��L�2���?x�����/��0�
S����pǎ�m>�7S����>|���k�G�u�-a6m�d�q�?K��9@��!�PhX��۵kgh(L�K;��yE�O��˼y�jV��\VV�V�mIv�/2C�rLX����v"������2oi>sʚ�g��Ί+췿����U::�����[�{5�j_�h;�i<��N`߾}�v�ڴ�F�����g�v[h΄��***\7����\����?O��{�Q�(�G��6��o~󛚶Y�_�m���}�ɚҡ��:�M�n���	-c@t�T��X�FtR��ׄ}��˴�VC��kE]�U+�@ԑ#G,,�����_�y	���hN�ڦ-[��[}:��<�����n���B1H, �(T�e���b۳g��E�=&, �$ڬ4�D��#�	Ӧ���`���9 �+���+�g��0m��	�!k֬�0��M��A|Ä�!�#4�*l�	l�P�B����cOB�_, `�W�La?��Hg�Ʀ��E�-[������
!˗/Ox?-P�s��hZ�k[���j� #`�	w���	���>B8F��ڴi��}��0,�5[�dI�	�*�ޠ�Q���1��Gp y, `;v������͛--Z�(�}�gY�N�,�T{M�S���壭[��[c�)�W\a �C�  �  �g,   �����i� �yN�U�*0-�/++K��0���T� Q�T��-���he�VA&�����c�������r�������{����Z��|Լy��)//�0Ӧֺ���0Y[�l1 �!`  ���������0m �*��<� ��h�E�� �K��lQ�B���$�ϼ�(���n�����_3��9�˱x�b�={����>o�дi��K_����ٳfމ�zٽ{�=���������*jx���ĉ�����륥��g����; �������[n�ŵͭ[�v�Sۼ�~����?lHΔ)Sl�̙֫W��s�ª6���wޱ(#`�K�.6dȐ:��Pad�������ݻ���`8�z���c�jH`�p%����2: ��s��6t��:�S۬6K��D��X����*7
��(C�l=g}��i�3uP�:  yB�J#��v��Я�EY�j�=��C�`�  1o�S=K���0h�p%�(J�7^�ϊ�����"=��1�+��ҤБ#G����8�߸v�ڴ�[�n��Y�j�,]���}�)  �i�J�ԋ��:x�qn5j�;l۶-�s�z�j�:��6o�\�
L��߫{9(j�F.ȟ Zj��Z�r�!=
����b#`  ��� @�i�ƤI��+աRݎ;��?�;+� ����W�,Y����X   >#`  ���  �3  ��X   >#`  ���  �3  ��X   >#`  ���  �3  ��X   >#`  ���  �3  ��X   >#`  ���  �3  ��X   >#`  ���  �3  ��X   >#`  ���  �3  ��X   >#`  ���  �3  ��X   >#`  ���  �3  ��X   >#`  �����lUUUv���_?z�������Zǎ�w��VRR�����o��y̯�7�v���{+**��K���������رcVVV�k�ڵ�؁��l}��>3 �K�-l�ȑ�gϞ��Q{z�ĉ�_1b��z�6�ȑ#VYY�kݻwwm���X��5�&&j�KKK�G��~�x���x�#`��Ç���Xt0�X]�tq�Ŏ;�>��x���ѣ�U�Vq����8n�:t�k�5&:X�,52�F���[����j,X �ԲeK���n�:�}:7��3ƶm��mڻwo�6�o߾ֳgOw��~fcK?�����u�'����������   |��գG�ꪫ2z�|]M�wK�z�j�z~N9�:?K�5�~�i����A�b~�m۶n�M�u�t��9��V����^uik�/��y����~������uk�g�z�����6l���:�yS��Օ�wӰA��%��ٳgE�]vY��r":��vV�ڜt{��[_�'���Н���߷k׮q{�ԃ�v-ި�z�4KAA��~���~w��x�F��{�<ѧO��ϫFR.�䒚���v������N���i֬�kc�����fb��d���	X��M�4������I߻y�w�<�a)�n�O��nV�2��|�;\���K�������wS��z7}��զ�͟����ü@���R˻�M'����q��6^X��U�P��eٲe��t�\TTT��Ν;m׮]�����m�v�v;�]�ƺ�Յ=+��8q�{_WA��[�A�?�>��^������6m����[D��ɓ��cG=�^{�'�T�[���hC�6m\�۫W/�q&�K~�D�R������kl� �	�T^�5W�}��,D�^����L�F��*��י�ք	l��Ŗ"���]�W)7��!�ޕ�h��Jnlڴɀ(�\�!C���[��E�7E�s�!`e����~�����d<M�N4qY݋�Λ�R\?�Nib�z@PW�� EN۷oo~�k��0�7yS�����/��zȀ(���k���M^V�??�>�@�[Г����3�h�9AB�ˏ����b�ڼ9{��u�ט^Z0��g.�V�}��?�S�N)}����1]~,����S�o�c���'5L�Ǐw�W�Νk@:�Rms��.]~_:9g�M���l?��BS��� 9S�N�Y�f�ڵk	X �!  ��X   >#`������@��U̲1zU�fOK A"`�3�<���Z�8p�]t�E)?ַ�������X B�7ިӃ�=��  � ԡ]2�]�y��9, D�g���JT��9K�Τ�Y��~����������0 �=es�NRب���w�"Qa�|F���$������ ���E��n��ݐ�:�m�f���/2~�6 D@���  },   �� �B�ɲ{�챷�z�ճ1b�6,������V��}��ّ#G �D�J�~��[�8�|wS �֭�u���M|��2w�>{��ޮ];��@^PhR�� ��������o�g�}֖-[f E, �ܹs]i��C�����]x�n����7 �* g����&
H��������Ν;��?��Ǐ7�>UҾ��ݦ˵'�Ǻoԩ���^�zYEE��^�ڎ;f �@��z����?n����6�{�6g���V�}�;߱�����&���������O>�Ģd���6q�D�\(����{uz���:��WPPP�9}�����~���@�!`���p���[�V�|�G������v��![�f�=��6t�P�5��S��b��su�]w�y�W�󥥥�O��O��G�-��b��ַ|�V4�k�;w�_��W � Ԙ5kVM�Z�b�-^��ՙ<x�]p�.�z�VVVV��,Yb���o"�<��~{�p%���.4�p�v�M7��mڴ�=�zNdӦMs��5�\c�������@�ਇj	����~�A����}�Q5j��XCZڳ�瞳��s6s�L�~qq�=��#�}�v�۷������2�~�ӟZ����g�������y\5<�M��8, � 8
N͚5s��5�W��͛����~����|0��J�<�L7�_EO�����+QP���/��B��Z���v��h��p�4@� `p�v����ڵ�*++c�gݺu5�S��d�(Ly�ʣE,���>�6n���E�3�w�� � 8�>~�{��'
���О��E,���.��P	�֭[�ѣG@�� �Q+j7���U����|c��v���Z/  ��X �Py�d�E��D�4��ǣyI%%% QD�P�&n��l�>����>ZG�U, ��׾�5w��_���� G[�4��-U�� QE��lݺ�ݐ�U�V��
~Q�R ��� i����n P��h3f̰�^{�N�w ��������ꪫlʔ)nO���� D@Z�&M��z��?�|k۶�!�nݺ�[EE�����>3 ��� %ݻww%fΜi����󵲲2{��7�W^��˗�J�Y���o۠A�j>�:a�ӟ��Ge�! �� $ԪU+�>}�}�K_��N;���ys�εg�}�.\��>}�؋/������X���:�5kV��w���d;v�}���g!�GX �5j�U�\r��|^B/[����?lk׮���<y�{�͜�̙�>EEE���}��c������vCg�q�u���������2 ����)gi��ȑ#�|m���nu�s�=��_�`�E���͛��TŢ
�͛7w難�����\�|�~�+_!`y���:t���j���3�x�{��mŊ��J�uꝒ?�0��5�z�y��U%��{�3��~�կ~e<��0����g۷o7 �G	��:ujM�<�ŋ۟��g7��ȑ#���v�����H��cǎ����z˪���G��C��}��6d��'X X�r�=��Ӯ������������3���xé
�{����[�N�@~ `p8��'L��n*��9W��Ҿ{��ĉn���RŪZ?nܸ��?�䓸���YT�@~ `p�>��7���_���1���\{��V\\l�������s�N��9T�;��������U�^�l��l<^ϕ�
�����n��n�G�v%.��b��P+�4	������7�ꫯZԩ܂��O>�z�<
W�{�v���qC=`��.W � Ĥ!-���^;��sݖ8
Z�	�y�۵~�z�ڶ/:UU��}�ڿ�ۿ�����V�~؏���i�{<*2���Յ7n4 ����Q��EÇ�����.��R���+kz]��;�t�4ko��s�&��k׮�{r�
Ƞ&�<��o��ܟu�Y�V��]�6HE\E�a�ji�P,�Kw#Y5�٤�J:W�^!B$/,ϵ6EV��t�o̥y9�y��l�����/|��j��C�6m�<"'�M�ʵ5��m��~`ӄpB�6m���ٳ�X�(`i��~��۶m�o���q�v�]w�9���k�W�����'q�W[�(��Vl�
���'z�gS:�G����{Bb�<�z������7�6W�2�uA���'J�Hӑ퀥�a:[�h����ڵ��R��C���AӉJCh�P�Kc�Ϛ��a����������S�.]����Z�w�g&�^���|(oN�6XVC���~���ĉݖ7ZQXYY�R�Vcj��򗿸�U�5W80�3�hU��[��,���=�HN:=Ӫ��3�mB��!z=<xЗ�#@��E��"馉���[�(P閊E����C���X�w�}n���� @�� �Ns5��� aD��h΂榤B!J�_4q<������6�@�9~�� ��X ��ʿt����J�?��mذ����[o�Y�*-���v(ݷo��/, S��"T��{��m��iE�׿�u��+����]M- �����
8MPO��N���6�<x�[�����՜�;w���߅^X����#��Bc{�Ţ�ѯ��s��I��N5zT�]u���i�_���v�7�%� ���m���SO=��ThPU�y���:���w�iP�P��?��?)?�_U��;�սӰ���Q���n�ͅS ����K�,��o��UzW�
o~��G�=~��JT/��R���G��z�T�@�� �F=`�SO�Ǐ�k��W/���}���wC���y�� �X |�~�z��eS�h5j��GX |UUU��j3f$���?, ��6Y-//7$�k׮�mEE��, �i޼�[M(۶m3$֫W/�߿�{�֭ ?� ����weTaѢE�ƩT����Dii��[�� ����p��ѣ�ꫯ��6��wߵ�۷bӊA��)���<��S�@��X �3f�7�񍔾G�J��֣M���_Z��I��R���z��{�Y�j�� � 8*r���X�|��q��w�^�����s����^{�~�_رc�@� `pTA|ǎ)}OYYY�ܡ����ҥK-JJJJRz�T�^�+����j�F�����/��w�=�� �G�  �  �g,   ��   |�����V�X���z��M�ĉi�~��ȶ���שӕ��ǏД6m�d{��I�{�^�%KՍӭp���\��a�r�a���mn(  @��   |F�  �  �g,   ��   |F�  �  �g,   ��   |F�򑶖ؿZ߻o�>�ѣ�5k�̐�ѣG���<��+((0 �}j>����8r䈵m�֐��DM��v��A�ر�5o�ܢ��哪�*۰a�;��c���VZZj���-[�+))�������U�ȶ[�n6`� -R;w�]�v���
W�W��~���[ħ�m���������t�:X��|�P�v�ڌw�֋p͚56|�pkݺ��!])\�*���mذa�, dv��a�w���1Ԇl۶͎;��s��C�e�8�xyݺu.dZT�2��ƍ3W�zA�9�Z���S��:�lْq��hxAWfC�1 ��L�Um{��qmm�^�umݺ5�p�Q���VQ����!�:��I=+
�����f:Â�Ѱ�޽{& B@�Uj���F��;Dl�1
V�λ��Ycƌ�Ĝ,Vt�W�
�N�eee֩S'�Ƀ]=NA�pC�Ν���8��5��7���[3j�(���t�%���m���-��2����`,z�N��J�6e�b���� �����Em��ţ���dhռ�d������� _����,%>)��Zw�>}�zr�N�~OǨOr���_s]c�ck�RϞ=-��2�UAS/Y��VM��gh�9@n�F{���_h�S[,U:��� O���
�0S��l `�+���P�N;��6W!.��,+MZ�d�'!.�9ϭ�l4� ������9�,ρ澪m��yX�4�]. �l��\���Z�@n�����f�V�K�B��rJV~N���T�5�l���9�����4�d��㠓>��-kW8<�@��V;в%�������mn~�uҋC���^mѮ];��l���rW�ځ���qρj�I��҃��:v�x��ψ:��o�>��
�XA�,�:!9'S��,���_�{��3�+]�vl�Q�)��O�ҥK�K�s����-���9(jg`�bSA3�ՄQx�9�d@W;J�AU��͚QY\f�uPP+����t���w�n8٣���i��z$�+C����իW�>ٽU�V�����i+�m۶������A �餬�m��7��J���G[�]P�-*���2�^�޽{����8h� �ztu���~��|�� ��������ҋ]���<�n�:_;t���-�z�(���������������m�ڵ�l�� ;t�P&�!���:n��1e@�C�a:F
B:mٲŗ���G�F�'zꄽw�޴C�G�����Çۆ2���!X5��f �G�hĈ�~���&b+@袍т�t>ҹ���8����>F)��|��^<���<!���8�'�+X5��7oNk«��4w��+ ��F��z�RݜX�zR4�Ќ����f��Ng���Y��]"�B���t�ze��J��6mڤ�}�$[TTd �O[��M5`u���-�A��-������"`���  ;ho�'[G�"  ��X   >#`  ���  �3��4yR�Z<-�M��V�+ ��[I��� uz�S�����Qū�g*0v�XC�T���Y�h�v.Ȏ1c��G�  �  �g,   ��   |F�  �  �g,   ����Ey7y �*��>��  �B��駟  ZX@�����!`#`@��}���N��mڴ1 *Z����
r\˖--����+O4��k׮DE۶mhJ�ڵ�\��   �X@��� �C�F���ɕ6���U� �='N��\���СCVRRb@Sٴi�Q�z�jkݺ�M����rA���G�ڑ#Gh*|D�.(F�a@S�   OE.`i>L��ۦԬY3C0��Rl8�����B�� 5o�<'��G�,���5k�Xԩ�x�Ν9����G���������-�Tp��i��ԩS��-r'UUUYYY�  Xt!�U�V�h `E��Ç]��?  8&=p��u�֍-�""�k�رv���

�W�^u��駟�S�,=w�СC����9���7(�>������7�h:tp�4�A��޽{��Y��Νw�����벴�Խ?o�<[�bE�G��ÚK�m��MF��L�L����M�M�K����K���V�a ,4wӻ S��9���;�8-��BV����\��ϭ^��粵!y���I�
Y�8Q �FV�������VQT��ɵmTԛ�+P]Y6� ��]�v��
���7%����;�5���F������]��t�����ڷoo �Q-��>���/��>}�!6Va��4ߎ"� ꣽ�m�X   >#`  ���  ���U�Vٖ-[��ZW�`���v�m4}ꩧ�|N�G���_�>�=�XMi�r�_oh	ֳgO��
7k;��***�^Ģڏ����'�{�basM45� ��7y������JAS�EmIIIS��a��a�=j>V��t$KW�Ç���رc�q�Ɣ����שq�u�V�,7�{�R��o��TL�<�NA�� dJme�^�5k֤��z�t�R�q:5�TK[y���7:�������b�ʕ�vBĢ�g���5��ٶm�!5�SXXX'�hyq�Kâ�CW:K5��w�^��rJ5`�љ8qb���֭K+`�7�N�ŋ3� c���o�ڨT�:�"{QQQ��j'SX�N�v���t�ȑ#�yģ�'Հ�v�v�������H+���N ��v!<��#`5]�h���WJ����c]���V7:R}�X�өS��`��LfKm_S����}������z��=X���ر�@m�1bD��c��m��5��;^�`�C������Q�Z�1�q2��������E�0��S�������#`5�`�L���~zQ�Hj�D�iӦY�F�]�c�
]����K/��  Y�|����S�f��t]{�0
\��m�B��pf2�9�˔�QuCjXH��蠧� ��^5��)d��Bn"`!#�-�.vvT�`iJ�BV��c�=,d�����d�k��  ���t!�I�'��1|�%�:�k�_��f���Ǐׄ,ڛ�բ:g6/Ǎ3F�'>6�;ਫ਼_��ɓg?��?1 N?��V�a������\�$d�5u������?�n�ߣ���ˋ-���w�cvy!KˢqR�*��8<�:u*3d�J�� ������k�����|GS��W�b�Y��� �O{����5�]��G���j/'N�f  5ڷPY���A� ��,���%��X�Ҁ�����͘�4h��:��b����X*%�l ��b"��>`~~�ȑC`���*��7�s����n�>��s�܀T?��V�)7�UUUu�r��U�ZɈ��    IEND�B`�PK
     �;\�	�2�9  �9  /   images/5119bd54-fe8a-4b53-af25-af94989a1f77.png�PNG

   IHDR   d   �   �R)   	pHYs  \F  \F�CA  9lIDATx���w�lYU?���d�aH�đ�DQ��CP�����A(
���)��/� T%���RQ%
�(Y�&��0$��h��o�{�>�O����}�����}��g��^y�}`�&\��ןu�Q��b���O�]�+��rr�v����}�&�{�d�����^z��K.Y�β�����E]�}n��N�娭�{L�����F��6A
ؗO���&���wF!\�Zך8p`�~mA�w������5���V�t�9�L6�~��Ǉ!�`�5l� 3K�C��l��ہ�����>zr��]m�c�4ܿ
�x≓c�9f�mk�M���_��F����������N2ގAdK��J��;�-D���V�	� }��� ;	;J0F���N��:m�igS�Zv� G`58B�=G��`�	B1�����Wmk�vvv� LIVR�1䥯����/nZb�
�
AJ��j��&��-��lR�J�ht��<e�X�t�Z�/�~,���K�+3Rx̫@��n;{vM�o1{ɫ��[YG`�d���	B?H��p'6N�Py�AV�Y�*��g�ђ�?dT���.w��r�)��}�s�s�=��D�эn4��-nх{>����H���w^��.�����v�<�f	���������'g�u�����A̎k\�������|���|���]7{��*�V���3�������_�~��|!�}(�׿�������կ~���o�����7��c��:�_����S�\��� ��5Y����K.�����@��|W�u(EY�3�����w�w���y�k_�Y��צx]�� �o;��+;���;ܡ��S�v�U�k��48Iu��3��d�i������I|?B�"��GNnr��tz��o}k'K]T?J</ĴSn��{Y��7���7�AGz���@ұҼ�c�_y��S��o��˶Z�l
�yꩧv�E��?��?w�o��s���nw��O��Ot����������悔y@D5P@Ǽ���ì���Z�N>����P��L���(d�{R����[�{�A�{d$wcF��@y�T	M�w��M��t�~�{�3�ַ��=�gֱ���Y�
��z׻^�.c�0�G���n���,4��ﺚ�/�����W�ڽ��׽n�G������`�~�+_���7���A[�b6�|�_���
��������G>2O�u�ް�:�C?�C��T��y�K^�q��W�M�mD�d����o��ށ m���}�VKtf�u�s��-B��o ��BL_��/�r&�1�0Ri�/�� :k����g:o���������_��D�g=� ީs��K_�R�����{'$�����|Ϧ���oi!�xB�,O�̦�V���R�Cxs1���ۿ�5N���>�=8T�M�lG�#��pD� D�dF�~C���8��\�P�C6��(i��ڂ�(�M��~��xr�;ܡW���٘�N1��ӟ�t������A��n��:�ͯ}�k��N:i&!S��B~�~C�� �OfgM�g20B� �5Bǫޭ	��d���FGw���\���JJ�ϞF�u�z����)�~
g���LY��}ϳ�!��w�˴�i(�:��R������������=�� G���8�|c����7�>W$���xΎ^U��U���ן}϶��)b��W�W3���k�9�+x%!���q��n6z�[1�M*�����G�<���lJ��3��ԉh��f��f��Ƈ�����3��c�z������-��~&
����w�^����WG�@����k�>��?��K�Bc8(�h�w��̃䴌�Ȳ�!J�~@\�)����������MwD�'@9��Z`��k����%Z�f��8�wm�7N�>��Y�ΪZ�ǉ�<F�l���D��
<S3�@G�y��߿렛t���!c�:�p�p���O�߽�s�%��,H�,r�w܃@��pa
�#n�N>��꫁��ȳ��!Y��ܗ%la �ҎvW1 �z��g�g'zЃ���I��o��o�3Rt� .1�����Ե�:
9��s!!�b2+��yMD�L�0�&��]�����<뻶b�!���G��ML�j�}K�c���$H�O�����!�S��T�%�e3�?�1���|���#<���;K��D���pr8b�>�c\n����6<��"�*H7��t�3��q*3#�����]�<uxf8��G?��I6�#�� ],=�!O}L�]۱"���H�$���
y�K���&���	y�����	Ô�y�Y~紭
	�/��I�7��M#`�O~��<u� �|B�Aز�,S��C�ϴ�km�ϗ��>��k��������)�>���Gj��!(��?�ӝrqC,"����˿t�ڴ�~��O=K(N?��N��w���A�J�ͦ+�����ߝ�6cZ��&<���*u�`tz�X�g�������*@��<D�$���d��ZK���w�=�>�Os� ��4FՁ��+7�������ro���ݜ��c�� 8��I�bLa�Y�$�y���N��z����w/��:r���$,�E<����n����w��]W͘��N����r�ې��z�݄Ҕ���n���DRy�������3O�}�{_g�����!.�T}�葾��5��i��8�>�-[*%ٶ}9���NTa�DD�9�O��Bz�T��\C~�3������R� ��27�\��0b�Ӽ����1�R���
����H9���3hz�.�v��L��̩�,(�K����DC��.��cv듰
d=2T��߉~"��x���{�pɩ�Sah����Tx$�=�#;������K�p	��,�s��Y�Y�C@����!۩>��bz�6�83O��Y4R�����;��1	�.�(�쨳��KTE>#
�h ˅�cZ����b�3�T�C��,*b��|�-�5M'+� �L�Crd�^���"�M*u��B��B~��y3��s?"YI�������37A��J=��<AЇ<�!�?��?��C~4��\�:�dN=�#��̩��V�Ѭ(7��?��\�F�ZpR�w3{�R���G�D$/�������N)u�#�ڴ1�S+�}}�����7zE��<��-\�7!j�*uz��@'��>�\�XV����ȏtdr��|�;�FqwB�����"<=�B���I��Lwpo2�y^��5�rDH`�y�&��O��~���<�w���-��)���?���y?�$h&�	*�0�BB,%JQC��CgP�%Q�03Ŭp����&��1J=�����f1D��Ї>�詛©�(󾭗����Aև��!�����d}�� B̴�$^������uaO~��DD��DD�C���"Y}�u�=u�o
�XFŮO�p]�e�x�� ��.�:��i�٩��ݮ�����$B�K�0>�At�o��of�q������"�x��G�|�_�� 8��J�$ٌA��뱾��"+tہU=uO����� Qy7=�	�vsr�����&H��Yf;En�"�pp�`6�p�tsּ�7������}:�E�j0�!eӞz�!1*���h��+&"�x�dw�S�̢l��m�1��M0T�zj��������gw/ջ��{C'LG7�0��o:�N�%���(�:�D��)2�L1؄R̆(R��e��v`�R�e�`2z�J�"��aj��|��R�ދ�p6䚁�_���8z%���S�t�3��r���$�y��*���c���M?��,�R:*��(fvB��  �	i:��Z^VJIz�� �"�{����ـ��ն]��F�H cA8R��[Փ�lE�� ��n@�h���oy���Z�/D1[M����I�V�ŝ���p���mo{��=�q��{������2s�� �O=뺻��O}���v ��'L\�X�\�*
 �שׁ,��{� �,AE�M�y�R���?��?����G��5s���g(󾭗�R���D"�o<q�(L��1BʈB�4B�XU�1C )Kx��Fe���*���$"b"�s�!+�mf N<�e��N.icaq�̌r���&U��YRS'��zC\���JPՅr}K�����ab�MO���3)M$��[9uHDh��$�.��|Q3���XU��u2úPʵ�z��S�"�+��:Y�"��Sӑ�ʩ'��pG�ev��f҇�N��"N���gXc�d�z�������;"dK�4{YZ�
/��Ωg �}R�D��#6����^()o�0D��'a�iCdY�=���Nw�e2Y\o{�ۺ��)\7g��n�ٝV�~!�g�]68�̒�W"�!��'ej�16���*�:b!ܭo}��J�"[xl�pe��2��~?��)�� �#��
K:�+�Z��Z����69�#��-i�8~�g~��!�7Ld�1�I6�k��=����ha`�ʰJ*��l����X�.Y�x�k_�Y����jz����r��O����z=�V9����/�,��}�>�҄�˒���A���ɟ�y��<�CR�r�{�{��>�#�X�����Sߍ%m%�C�V����߳ <���8F]b�������Q�e޷��V��~��{�ʥ(#�����Uف-䐧N��&v�6�p�����:	���9�P~<ubȴ�4y껡��2D�mg$
O�3�����l�SGQ�����<��P�d�X"�k蛚Z|�ZCT�lg������|�o'!�IbW�YR�&A�Sw�\禬joݗmb/8�N}6�e��K��J�#\7C���>�D��ʯ��L����/��W����8S���������9$""�>s}�S�rφ�n�%^~D�_�'�aqJ]mt����S�����I*_��k�y괿ӭ��R_�ʀ�.�&"Ϙz�S����׽��:n�3ͺ�쁽߭B:�Կ�ԓ�h��2�g�z""tɂ�nVd�*����ˏ(��AK��m<W���:Ecf �c8�Q�WA����V�;O���/	���!��N�%<�l�߂U�:��j�V����ԉ7�Ea_""��Y�I��C�l�U��o����\���a~E���,��p����Ϙ��eJݟ]t��կ��tZ39�������� 7c/�G�s��'�bo:�Z�枋��Tb������͈������v������u'O��ES���}r�@���W�r����K�Tt`� �\l
�RfӂL��>��3���v��SI�^<�9�'�D�?�Q��y�-��M]�<�%5wU��򘔲�g5��)u���.�<���L��1Squ�䤓.�s�\�q(��S깏��Ĕ-cS��[��z���x̲��p')1��Λ��J=u[��F��˯7ڵ}�UT���&̼�۾TN�x�L��*�G�d�$�����J<�}�� �] ��7��,��R���!O�y�
�ó�<u�#�W��
�V�q��m9����L��p�7^ �zի��ƟUR5�-�-���MtC�A�A]�Av�ɟ����	�Ѓ�!�O]鏙�:�Z��S��S�R�A���u�JX�d���,?��
3ξ,��~�(9��S���C�e9���gq�� 9\2�����9sD��o��UA�B#-1Ԃ�W<#
+�����=SߜX��T�/��� {�����dÒk.;�e�~�9"TyR�q�^S�M���x)��.�"��;���Lc�Cr����ۻ,:���/�L:��3'�w�y���6��M��?��?����]!���fà$l�e����hw�_��_tVH�A�Y�Qd���_�W��wow�T�&.3�#�v��G��ɋ����̩�kk�-'x�9�I�s�e�@�,��PH�� �ʾ C�����8�a/������<�T��'�R}bR��_�x�ln.��9���:G�.�d�����ؼƿl��׼f�h+��,t���k)�.�jA��6�Q4ۘ��wQ�]��pн[_�x�b]�ԍs� .����x�DИ��Z@�w��1���d��M_��u�KG_���?�a�l��)�\���g��S�����!�+�e!	O=;{����0�ť�PB�:do�e�AN���������i���)��+�$�n3[p%q�!�,@��mby�p�of����<������^C�z��^}2��� r��79�?��?���ǿ@I��^"*Q��41������)��s�:����ΞfƐ����R��_�=���L�>���������ʃ��3��]�"�J��3�pYG\��N���Їv�/|��"9YYx���M0ق��\o���l��YJ��c�ON<��_|���2���[�}	���3���/�RW+��W���~e7�ܛչL�*k�� !�CDL%N}��q��U|����ٳ!��驓�q�s���˯���ך��7�\r��/�����?|�d_5����|�:
cd?���&Y-�� :�>a�հ���g��㝢�V=',����9V栧.4lJ{��\ȁ�&��&_<�;�[��^$_u����3x�w��Xz�����l���K$����p�~��X���J>�F��	n���!ӣl�d�nu�����&��<�~�eK�t�/�e�B$A�ѱ��+ׁ>�W��WӖm5�3V#�hvl^�B���`���&���9�����4�9�~w[�}���3�:���.a>g�
ʤX+A�)(��7�[1J+��93�	��Ѐ��^�Գ7HQ�-����[u�l�t2�T�CC����>�)O�Jf���7t����S������W9�y(��z6��b'�Y��7J��e�&�%�H�7�:�O��eoy�[zO�IU|��~�Ɵ�>�e���F�P̘�S�ᡘ�,?�a96(c)�8��l�'	ߔ}6������[��kD��2vN��vO��M+�1;�ό�Ⱦ]=��X���x���d@��W#'fG�$;B佁4��̂��3�:<��S� ϶����qp%�q
� g�\������/KYl䮙h�Me
�.��Y�[i���sω�,x���,C(=�1;�� ���>ީ4)�#���!t�|����{o<ux�C�s<ubAN��O=�� �b�>��O�)B�Zs(���bc�����O=���f���	vB�����,�Fə;Y�	�o�������B�=�+x���Y��ڤE�U��c*̂�1P�	忽B��S�?(y��B
7��	�F��X�M��PC:C? ߌ���y�����|��!	�mғ_F�(�ҁl���D,���m���1tA�D��SO�=vC�$������߾'�/Jj"��0
y�G�1�l�D�Cb߲�D̙�fA"���Rhm�`����d�hI�n@�x��rDEy�!�$��g8�f�~Yq�X���胤�q�>��k�J��q��SO�Dj�|3 ��������su-W-"\�8Ž6��~v�K���e-)� }~����p�8&�<ԜI��M֩{�.a��v� 5�LI?ŉ��ܕ9t��M��O���u�`	ٹ�;�-x�Y��͌0�g�5���Di��=X0�q�<����NL�<^)�^�ԧ����f��f+k�S'�x��&D�K�:H��P�(E���La,�j�V/�Po�}6Y��ԍמ@c�Sgߛ-�"��7}���J�:�Ar�Μ���n:!�^��$R�'�SݯR�RO1ɂ��D���D�nƌ-ӿ �ܽ,J����-+����J�Z�!�v2e;7��r��I�rb���8�� �&Q�����U~:��Y�;��<5Y�ԕԳ�6uN�*��oGg8(�@"F$n�W	���_��_7��p�c+*b&1���ʀP�������ߤI����3$������}�.E{���ED�9�M2���s3$G�r��n@2k�����ɽll��v%�ʗ����LJ�x���M3b�2
���MO��ޣ�/Ο�@����sN*%	̐O=U٪�y�<H�⩗����NE1���������N�E��˓�`�"�)щMO=e��*�J/0�R��%h�;��ۿ��p����눓G���"�������J_���E9�g�?��4���֔;���(WB,�'>��
'�G{H�W��՝�D��ٟ�٬b�	OxB�.ɤ�R��`�	TE����wr2MKυ`��w�sq�U���Ru������I�,�S�h!l�C�P�X�)}m.G�����:���g�uV�	 B��R^:�0��"U����s  $ty�-���ĩ�D+���$��pih�6+����L�sq��se��!H�py�WvBr���gǈƔ�JHN'N��tu�*r��:۽"��
�MvN���j]�H���3���!^-��_�����`9�ק�Ax���om���Hym��K>�OC� �F?���Bb�{[�׳�a�܊w!��9��þ�b��u�Uw[���zy�HA�����ǖ�++O��M~~��%K���HYi���2o�Bj�̿���\����7�q�pɔ�d��N��G�������)N�������kv�ip��Q�i\���25������.b@ܖ��,9������=�3.��S�̕�S��Xt���9b�������NV�6�_���82Gݕٷ�D���ĹrȌ�s#���	q��1vGHP�DorD� ���t%�1��jv�p��ݯӛ��ǘ�Is��'�Q��0CJ�k�:a90X'�-,��l�=�gg�G:{�[ݪ�b(rB9sP3��vޛ3�p;�k�G���������Ɋ�0��x^|(�1!�'�?�DJh�ya#�x�L��1G�Oj.�9��X�阍�Ӊ���)%665q�
A�P����`�Rk������=��� c*q~wDĔ 9`�'ֆ�xY(Q�	���L$��!}�v�a8`�ri`<uYYˎrb��zr�����z���!�0���rݿl��n":�u�gjF)By����GT������	�Ր؝~�˒�{��(�a�L�5P�K�?�B?چ�x��c��O�@D��ڊI�$D?�!�LE/(�.'��ܜ��A�uS�W[*Y���Y�f�X}��lF��`Dd�1���w�
���1N[2!��:u <l�"��'1��zj��i`�S�����<acG9����4�{�'�⓬��֥��DT�qG��3R>�7v�? gD1Q�=F@�r	(zy�?*!֏N�����X	�͒��ps��S|s�1��ίw����F��p�}�s;/Db��>����0 �� �]v�9Lě�w�'a�q�91�;��N�3ͽљ�YֽP(W���du�5d�"bQL����:O�_:�<f+ǒ���s��x��ǃk�N�,��A
t��8V9<v��>3Rʱ��7���j7Fk�~� �@��}�\�cE�M��'F5����"� �x�1\��< '��7������!jz_�4x2�%��Z~v�;�>��7/2�60%�����ߓ�.7�Y�eƳ���"0Fw�㖼73ap�w�?D��߮�
��ʀ�ffq��q���ˬX�As��WP%������AX3�ٓ�.�?�\38\s饗L�=F�|��yW���-��/���Go�Q�P�c -jtߟ��vc�[�O3�g��q�l�8��@��;<��҃t3p��p�fiЋ�N"��Ό�6��;[ۀ܋��>�}�\Kdy��lDGQ@gb"\��bl�f�;AL���Q��cd+)���g'��y�S��z�Zv{	.�+�<�n���	qw��fPL䬇C�Xl�~����5��?��]�C��d�w$$��,�b�%~W����iE�"��<��iA��W���;�n����C/e]q�r�q:d6���Dݡl���D�5 �f�F�����~
�s��Q��DK�y�O�6�1
]�!\��E -�����x��C�ܦ�.8V�/B��\�˳H1{� ��"�kzv��,)�%�ͻ|� ��|w-˦˰���"��tv}�q�����O��a�$�Ce�<3`��z\�d�(�riV%���A�2j[�\cʌa��cVP2ٴ&'�x?�ā�u���)H���٬�;D�>����A�lh�)�s�M|�r� ���MO=���_��n:	E����(S�!"�C��^�I�;!��0��Y,�	I���14�!޸|""Q�&vVu*��W�'��g_�����E��ݍ,.q�:ܝ%���7M� ٻ�M�[�7�,�����������D{�^G�@,&�����+uk zNi���C�P��� ;�9vT�d�� \L�e�Rb[�{��Y��Z�+�{)��D]Jl����ȧ�͒��l����kc��?�e�b���eVJ�A��~3���r�8I�N����[[q����@��ُ�a ���i)���k�����1�����l�Nt���	[D�H�+��v��-��(�>p�0>1J%p�g��=�Y9�8YR��	� �K�Af^ć�Q��&����!��Ϙ�"��)�t���uM}�c�e�Lɜ�����)y�x���9O�P0n��|ñۭdٰ�:�2��٘��Ѿ��NC�Q̒3Əa0+����(y�x�l��{�~l�L3r�8����9U����eiN�X�k�˾���B�"f���E	I��=~g�E���2���������:�� K��J�t��ZHLX����!0�����w �2����z-�븴�(�������&g%��x����YG�y7�qj�D�#��c����3q5詧*�׉���:���d�g�SqB�T�5Q���{R�h���� �)��}�R���k��k]H�y�{�,�I4:���Sf.s	y�(q����Y�i�tə�׷�L"�NiCI�^O��b�∱Kٲ�.�9�5~ғ�ԵW����
��M��c��m�/���ݟ��gw�2�]*�2��1��1P�Q����g<��OP��#R.ݪ�9z��˷
����`�^���62�v�}Y	Ь~�R��b9��Cc��h+k�P��/��?��w&�|���g?��K���?ar���}`+_m� �<�6��׽�u�S�k�eS�������LVO	j6��o�V7Cb�v<m[������O��c�ȻrKd�����j�����k'��$~�AKQ�ʚ讱�����t����9WM%���}wr�'?1��mo7{�������ߚ��U�\����h6i��8��g?3���R��n�L�Ɨ?��ɩ���d�V�CV]�8�繖R�M��ح�p�'G�^QeƯ�j?_�q�i���%���v��)w^0�'N�{���\f�O����ɿR1_����0{/�1ځ�'Go͆n�H7L�w�7�1���o0˺;%�x.k�D��Egc_��2����8�P�u6}��;��q�)�1�\�h��,�z'��Η�Df}K	��bc������e3� Q9&�}ܱ�+Ubԝ���\H�oRz�"�A��J����ʦ�;���M�ۻ�ҷ��.�;�&��.J� ��{2sCк��1f�	L?�?���;rq�C���)1�/��L�8n�A�S��s�e�?�|0�df� ��T�O�8����-�4!�Ut�w�T�+&�"f��l�e���
�M��lA�t ל��S]r�V�	Sy}���|e7�+g���L�n�����︆��l��z�T\�<5��m͑L!g��$W�_]fZ�=�S42z$��Tr�
���,�Y��6�S ��ܲ��Ny�J|>�9�Y�C6t�w�C���y�?'���Xs!��/��ԧ>�[O����I�㈬ٲ�ܘ��J1�"�E*c��-E�{��b�L��}�B��w3)����u��N���B�V�*WU�O=��b��KԈ(8zֳ���g��՞z֩s�<�,I)'s��d���� Pl�S�X��e�'�`$B�_ȓ��бہ�Br�)R�;�Yn-�����?�ѿut\�& {�x7���"�k�%�<2��u��3=�l+kXޓ���}H̀ٲJ���X�sWI_��EY3@�d���*O��-�݂�8m�Q"����:��5B�1I�><�����q)X5��>�D6�����B�6b��/�dp���_�C�L�X�-�"�[��lLdH�JU��B
��)+@��y���ڊ��̤kŁD#:WoH ��$�t�7ҙ�.k��e�>��lnQ��:�����5��<'��j-i�4�,�����zG��iO ��	Z�M�����'��{������cd�ex^�:���;�9C��^/_�]Ct�Pۮ����5��Wt��r��%��� !q�pV`\�m-~��ֶl
��/��!e��T~�S��V�rS=Yߗ�O(����d�Y��jU���\���U�M����g��B:,�g	k�76uYr_]�Q�N��0�!=�L�P*�k2$����-A���!��kUZ�uq���W�Z�	*�MceB-$'����Ͳ&��d��[K�[Zf�Fqu2�˜�,�چ�uf��d�|K�ؠ�D�Z��x1P�a��E @�KbMX�׭.�>C�ʗ~���:m-����Y�b���#0�h�*���-�����EɫǺHu�^�owDZc ili�$�R�:�\kdR뎬ұ�c�ۊ.��|{���38B�=G��`A�냲�61�2t]������v�G�]+7�,������Ӿq.%Hvд�,9�$oR��AK��w68$�+�I~�Ɇg&��fݹ�t�2Y�����f� �q�&�����RKl,|"x2N�f�l�q��i�bK	�e�A���s�kK���h��鬁pƿYg�\#��v�D�[@�a�l	�<Ū�̳�(}��b�6N�>��Sg{�,�O�EQ�x�f�
K!��q%� -'�/4#��2�t8eE���Y���H�oYL)Y=1��K[�����U7�цY]�d��\_e�q�W���9Z���VD/�����
��������q��Ii��5�����0D��8U�D?�:N�"�h��O�n+�XN�U rt�g!V<(�¬	}+�0k��(X�R"���;Ye��u���g�e�n�nk�gAdK('��^p6 Q���������}_�Z}]X��C������!ʿޤ�7�z/uf����Ap�+_���~��m-��D�휊f���N�͛�A���}�u��g�<��C�ғ���Dn
(�f�"JU͗�cVYsR��r���u�8[�g��8{	�&�t6ì̢M�V�:�5e<u~�xaIi�܀��
  V�F�>�A$)��G���ԩ�I�Xk��^�q�m�n�e_k�q2��Uz�8]+��7	�U�o����͒�\���1\�Q�!���#˽��ö;��zcJ��=�W_���'w�2��yQ%i�"��z{%HvM�d��q���E8��/��ϲ7��11F�q��,U�`Pd�2�e&�SnU���s ��	1�@&�.�#9d�`��`�E�0�ȪgB�4}�����G}�[J�e9��@��>0��`�>��Rd���:�u`'�8:�e�	&n�_�k��xѭ�����C���W�P~�8�5�M���WrOf[T0�����ie��I��az��Ob����]���:X��v���48C#Q	���-9�Pv�7JX��1� �qֱ�M��
�b��2{�:�hm��my���=�90���z#��]�7N�`�ғ.�(c�ɰ�b'�qanĲq��r������L�1���R��0�fL=50[�
��*R=� �͢U����ٵk{ׁ��
u_W�����ѰxR���c7�C�@.��f�fK���7b�^��Ac����#ډ��d-��s|D��7�Y!��
[lj��MB�G�@�����Y��3a<�����`�ho2�)N:k�:����K�K���*c�U«�3a ��5�>M�Q�!«B��U{M|�u'�E��g}k1jہ����J?��n�s)A�}d���E�� �/��%#ȼ<�!�@�\u�e�`Z��za�\�C�}�Bj
A���i���kwx��E9k�Y��lv0�Xh��B�r��ԓū.!��2Βh1l��b��4�lY�SL������{��f�{�V��@lP��eG%8ּ�$0�YC9��'����o� C9�@4����Ӗ)<�14�{hY��Zr ���SƘ��)^�`p<U�%��f�>Ӫ�K^�n��պ`�/zы�B<K�j�/��Ƅ)�-����w'�m%��S��f���0��uv��˦���ĹU��s�B��A������6�|�j�5[��=SG�+�r5y.����q�V��/��Bߝ����~������Ic���i�������΍�����u�B��O?�w�>��gLe�k�	W������3���g��;S��'&�q��~�Td�`ڏu�y���+��k[�ή�y�c�;�i��긄��$_čB�$    IEND�B`�PK
     �;\�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     �;\��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     �;\�	V���  ��                   cirkitFile.jsonPK 
     �;\                        �  jsons/PK 
     �;\>�a)  a)               3�  jsons/user_defined.jsonPK 
     �;\                        � images/PK 
     �;\<jݍ�� �� /             � images/f679dfe1-7b61-46f4-bc7c-d69b61239140.pngPK 
     �;\ŏjY�-  �-  /             Ǿ images/f78ae6cb-3b21-49f8-a0a0-4b83f9561715.pngPK 
     �;\;+z +z /             �� images/47e6ec23-9fd2-4f79-b93f-ab3ba2a25103.pngPK 
     �;\�	�2�9  �9  /             !g images/5119bd54-fe8a-4b53-af25-af94989a1f77.pngPK 
     �;\�c��f  �f  /             (� images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     �;\��EM  M  /             V images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK    
 
   �   